SV	SN	chr_1	pos_1	flag_1	chr_2	pos_2	flag_2	qual	sg	calling_type	simple
C1k_FP1705220210LD01_1:1060743:+_1:1061672:-	FP1705220210LD01	1	1060743	+	1	1061672	-	14	somatic	DSCRD	1.0
C100k_FP1705220210LD01_1:1910926:-_1:1963488:+	FP1705220210LD01	1	1910926	-	1	1963488	+	19	somatic	ASDIS	0.0
C1k_FP1705220210LD01_1:2840012:+_1:2840732:-	FP1705220210LD01	1	2840012	+	1	2840732	-	10	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_1:6331484:-_1:25787200:+	FP1705220210LD01	1	6331484	-	1	25787200	+	50	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_1:6387047:-_22:41740688:-	FP1705220210LD01	1	6387047	-	22	41740688	-	22	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_1:6387054:+_22:41739996:-	FP1705220210LD01	1	6387054	+	22	41739996	-	49	somatic	ASDIS	0.0
C1k_FP1705220210LD01_1:9490188:+_1:9490883:-	FP1705220210LD01	1	9490188	+	1	9490883	-	19	somatic	ASDIS	1.0
C1k_FP1705220210LD01_1:12706692:+_1:12706895:-	FP1705220210LD01	1	12706692	+	1	12706895	-	13	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_1:14029349:+_7:45483760:-	FP1705220210LD01	1	14029349	+	7	45483760	-	99	somatic	ASSMB	0.0
C1k_FP1705220210LD01_1:14954223:+_1:14955026:-	FP1705220210LD01	1	14954223	+	1	14955026	-	40	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_1:17861583:+_14:89079951:+	FP1705220210LD01	1	17861583	+	14	89079951	+	29	somatic	DSCRD	0.0
C1k_FP1705220210LD01_1:20244031:+_1:20244857:-	FP1705220210LD01	1	20244031	+	1	20244857	-	34	somatic	DSCRD	1.0
C1M_FP1705220210LD01_1:22086175:-_1:22755433:+	FP1705220210LD01	1	22086175	-	1	22755433	+	22	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_1:22157719:-_17:5278289:+	FP1705220210LD01	1	22157719	-	17	5278289	+	23	somatic	ASDIS	0.0
C1k_FP1705220210LD01_1:26467605:+_1:26468054:-	FP1705220210LD01	1	26467605	+	1	26468054	-	35	somatic	ASDIS	1.0
C1M_FP1705220210LD01_1:27030859:+_1:27180255:-	FP1705220210LD01	1	27030859	+	1	27180255	-	61	somatic	ASDIS	1.0
C100k_FP1705220210LD01_1:27335883:+_1:27355490:-	FP1705220210LD01	1	27335883	+	1	27355490	-	21	somatic	DSCRD	1.0
C5k_FP1705220210LD01_1:28865563:-_1:28866603:-	FP1705220210LD01	1	28865563	-	1	28866603	-	81	somatic	TSI_G	0.0
CBeyond1M_FP1705220210LD01_1:28866596:+_1:47542042:+	FP1705220210LD01	1	28866596	+	1	47542042	+	59	somatic	ASDIS	0.0
C5k_FP1705220210LD01_1:34981001:+_1:34983343:-	FP1705220210LD01	1	34981001	+	1	34983343	-	28	somatic	ASDIS	1.0
C100k_FP1705220210LD01_1:36882993:-_1:36924206:+	FP1705220210LD01	1	36882993	-	1	36924206	+	42	somatic	ASSMB	1.0
C100k_FP1705220210LD01_1:36935134:-_1:37030901:+	FP1705220210LD01	1	36935134	-	1	37030901	+	17	somatic	ASSMB	1.0
C5k_FP1705220210LD01_1:42243366:+_1:42244862:-	FP1705220210LD01	1	42243366	+	1	42244862	-	27	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_1:44560428:-_8:131711090:+	FP1705220210LD01	1	44560428	-	8	131711090	+	44	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_1:44561464:+_8:131711078:-	FP1705220210LD01	1	44561464	+	8	131711078	-	29	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_1:45244132:-_6:25744294:-	FP1705220210LD01	1	45244132	-	6	25744294	-	62	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_1:47021482:+_18:68889067:-	FP1705220210LD01	1	47021482	+	18	68889067	-	22	somatic	DSCRD	0.0
C100k_FP1705220210LD01_1:49067990:+_1:49079246:-	FP1705220210LD01	1	49067990	+	1	49079246	-	93	somatic	ASSMB	1.0
C100k_FP1705220210LD01_1:50179051:+_1:50227686:-	FP1705220210LD01	1	50179051	+	1	50227686	-	99	somatic	ASSMB	1.0
C10k_FP1705220210LD01_1:57552661:+_1:57561455:-	FP1705220210LD01	1	57552661	+	1	57561455	-	41	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_1:68585935:-_12:61567903:+	FP1705220210LD01	1	68585935	-	12	61567903	+	33	somatic	ASDIS	0.0
C10k_FP1705220210LD01_1:71086571:+_1:71092180:-	FP1705220210LD01	1	71086571	+	1	71092180	-	99	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_1:80599652:-_7:100016522:-	FP1705220210LD01	1	80599652	-	7	100016522	-	93	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_1:84360081:+_12:3608319:-	FP1705220210LD01	1	84360081	+	12	3608319	-	27	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_1:84899835:-_1:106063080:+	FP1705220210LD01	1	84899835	-	1	106063080	+	67	somatic	ASSMB	0.0
C1k_FP1705220210LD01_1:96598407:+_1:96598816:-	FP1705220210LD01	1	96598407	+	1	96598816	-	49	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_1:97450821:+_11:22699899:-	FP1705220210LD01	1	97450821	+	11	22699899	-	63	somatic	DSCRD	0.0
C10k_FP1705220210LD01_1:97530623:-_1:97535885:+	FP1705220210LD01	1	97530623	-	1	97535885	+	80	somatic	ASSMB	1.0
C100k_FP1705220210LD01_1:98948607:-_1:98987980:+	FP1705220210LD01	1	98948607	-	1	98987980	+	21	somatic	ASDIS	1.0
C1k_FP1705220210LD01_1:99551783:+_1:99552379:-	FP1705220210LD01	1	99551783	+	1	99552379	-	69	somatic	ASSMB	1.0
C5k_FP1705220210LD01_1:103504515:-_1:103507514:+	FP1705220210LD01	1	103504515	-	1	103507514	+	15	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_1:105563674:+_1:189721188:+	FP1705220210LD01	1	105563674	+	1	189721188	+	19	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_1:106508532:+_14:59221145:+	FP1705220210LD01	1	106508532	+	14	59221145	+	32	somatic	DSCRD	0.0
C1k_FP1705220210LD01_1:106787248:+_1:106787684:-	FP1705220210LD01	1	106787248	+	1	106787684	-	24	somatic	ASSMB	1.0
C5k_FP1705220210LD01_1:106979939:+_1:106981337:-	FP1705220210LD01	1	106979939	+	1	106981337	-	19	somatic	DSCRD	1.0
C100k_FP1705220210LD01_1:107187826:+_1:107232687:-	FP1705220210LD01	1	107187826	+	1	107232687	-	49	somatic	TSI_L	0.0
C1M_FP1705220210LD01_1:107213409:-_1:107451488:-	FP1705220210LD01	1	107213409	-	1	107451488	-	87	somatic	TSI_G	0.0
C1M_FP1705220210LD01_1:107217816:-_1:107477306:-	FP1705220210LD01	1	107217816	-	1	107477306	-	87	somatic	TSI_G	0.0
C1M_FP1705220210LD01_1:107219087:+_1:107524722:-	FP1705220210LD01	1	107219087	+	1	107524722	-	18	somatic	DSCRD	0.0
C1M_FP1705220210LD01_1:107219885:+_1:107445679:-	FP1705220210LD01	1	107219885	+	1	107445679	-	18	somatic	DSCRD	0.0
C1M_FP1705220210LD01_1:107228856:-_1:107916257:-	FP1705220210LD01	1	107228856	-	1	107916257	-	55	somatic	ASDIS	0.0
C1M_FP1705220210LD01_1:107234374:+_1:107405987:+	FP1705220210LD01	1	107234374	+	1	107405987	+	14	somatic	DSCRD	0.0
C1k_FP1705220210LD01_1:107285149:-_1:107285522:-	FP1705220210LD01	1	107285149	-	1	107285522	-	42	somatic	ASDIS	1.0
C1M_FP1705220210LD01_1:107285591:+_1:107721211:+	FP1705220210LD01	1	107285591	+	1	107721211	+	20	somatic	DSCRD	0.0
C1M_FP1705220210LD01_1:107287867:+_1:107572188:-	FP1705220210LD01	1	107287867	+	1	107572188	-	26	somatic	ASSMB	0.0
C1M_FP1705220210LD01_1:107297440:-_1:107717067:+	FP1705220210LD01	1	107297440	-	1	107717067	+	99	somatic	ASSMB	0.0
C1M_FP1705220210LD01_1:107400671:-_1:107910578:-	FP1705220210LD01	1	107400671	-	1	107910578	-	50	somatic	ASDIS	0.0
C1M_FP1705220210LD01_1:107445680:-_1:107635812:-	FP1705220210LD01	1	107445680	-	1	107635812	-	57	somatic	TSI_L	0.0
C1M_FP1705220210LD01_1:107446168:+_1:107551055:+	FP1705220210LD01	1	107446168	+	1	107551055	+	33	somatic	DSCRD	0.0
C1M_FP1705220210LD01_1:107452094:+_1:107635856:-	FP1705220210LD01	1	107452094	+	1	107635856	-	43	somatic	ASSMB	0.0
C10k_FP1705220210LD01_1:107477306:-_1:107482496:+	FP1705220210LD01	1	107477306	-	1	107482496	+	34	somatic	TSI_L	1.0
C1M_FP1705220210LD01_1:107511920:+_1:107694670:-	FP1705220210LD01	1	107511920	+	1	107694670	-	71	somatic	ASSMB	0.0
C5k_FP1705220210LD01_1:107544401:+_1:107548791:-	FP1705220210LD01	1	107544401	+	1	107548791	-	35	somatic	ASSMB	1.0
C1k_FP1705220210LD01_1:107549646:+_1:107550009:-	FP1705220210LD01	1	107549646	+	1	107550009	-	43	somatic	ASDIS	1.0
C1M_FP1705220210LD01_1:107577766:-_1:107698577:-	FP1705220210LD01	1	107577766	-	1	107698577	-	51	somatic	ASDIS	0.0
C1M_FP1705220210LD01_1:107579789:+_1:107698702:-	FP1705220210LD01	1	107579789	+	1	107698702	-	50	somatic	TSI_L	0.0
C100k_FP1705220210LD01_1:107579849:+_1:107649066:+	FP1705220210LD01	1	107579849	+	1	107649066	+	16	somatic	DSCRD	0.0
C1k_FP1705220210LD01_1:107661965:-_1:107662355:+	FP1705220210LD01	1	107661965	-	1	107662355	+	44	somatic	ASSMB	0.0
C100k_FP1705220210LD01_1:107662029:-_1:107679719:-	FP1705220210LD01	1	107662029	-	1	107679719	-	68	somatic	ASDIS	0.0
C1M_FP1705220210LD01_1:107663319:+_1:107916318:+	FP1705220210LD01	1	107663319	+	1	107916318	+	40	somatic	DSCRD	0.0
C100k_FP1705220210LD01_1:107695111:+_1:107713637:-	FP1705220210LD01	1	107695111	+	1	107713637	-	50	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_1:109078068:-_2:166174925:+	FP1705220210LD01	1	109078068	-	2	166174925	+	20	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_1:109079177:-_2:166174817:-	FP1705220210LD01	1	109079177	-	2	166174817	-	33	somatic	ASDIS	0.0
C1M_FP1705220210LD01_1:112965980:-_1:113209462:+	FP1705220210LD01	1	112965980	-	1	113209462	+	40	somatic	ASSMB	1.0
C1k_FP1705220210LD01_1:114436863:+_1:114437856:-	FP1705220210LD01	1	114436863	+	1	114437856	-	20	somatic	ASSMB	1.0
C5k_FP1705220210LD01_1:120366968:+_1:120371799:-	FP1705220210LD01	1	120366968	+	1	120371799	-	30	somatic	ASSMB	1.0
C1k_FP1705220210LD01_1:145694081:+_1:145694344:-	FP1705220210LD01	1	145694081	+	1	145694344	-	91	somatic	ASDIS	1.0
C10k_FP1705220210LD01_1:150022545:+_1:150027974:-	FP1705220210LD01	1	150022545	+	1	150027974	-	20	somatic	ASDIS	1.0
C1M_FP1705220210LD01_1:150392175:-_1:150568164:+	FP1705220210LD01	1	150392175	-	1	150568164	+	57	somatic	ASDIS	1.0
C1k_FP1705220210LD01_1:151037213:+_1:151037611:-	FP1705220210LD01	1	151037213	+	1	151037611	-	14	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_1:151278094:+_1:162538266:+	FP1705220210LD01	1	151278094	+	1	162538266	+	11	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_1:152610787:-_18:4218827:-	FP1705220210LD01	1	152610787	-	18	4218827	-	99	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_1:156407795:-_1:211022624:-	FP1705220210LD01	1	156407795	-	1	211022624	-	99	somatic	ASDIS	0.0
C5k_FP1705220210LD01_1:159020887:+_1:159024418:-	FP1705220210LD01	1	159020887	+	1	159024418	-	32	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_1:161930887:-_12:39860506:+	FP1705220210LD01	1	161930887	-	12	39860506	+	33	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_1:164277385:+_1:228881161:+	FP1705220210LD01	1	164277385	+	1	228881161	+	23	somatic	DSCRD	0.0
C5k_FP1705220210LD01_1:165428983:-_1:165430339:-	FP1705220210LD01	1	165428983	-	1	165430339	-	43	somatic	ASDIS	1.0
CBeyond1M_FP1705220210LD01_1:166723266:+_1:215556899:-	FP1705220210LD01	1	166723266	+	1	215556899	-	99	somatic	ASSMB	0.0
C100k_FP1705220210LD01_1:176116783:-_1:176131865:+	FP1705220210LD01	1	176116783	-	1	176131865	+	48	somatic	ASSMB	1.0
C1k_FP1705220210LD01_1:177082500:+_1:177083213:-	FP1705220210LD01	1	177082500	+	1	177083213	-	80	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_1:199500696:-_1:238615390:-	FP1705220210LD01	1	199500696	-	1	238615390	-	71	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_1:201783847:-_1:244309004:-	FP1705220210LD01	1	201783847	-	1	244309004	-	99	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_1:201970618:+_1:244584072:+	FP1705220210LD01	1	201970618	+	1	244584072	+	35	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_1:209132347:+_5:109480197:-	FP1705220210LD01	1	209132347	+	5	109480197	-	26	somatic	DSCRD	0.0
C5k_FP1705220210LD01_1:211021606:-_1:211024542:+	FP1705220210LD01	1	211021606	-	1	211024542	+	91	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_1:217404493:-_3:158848652:+	FP1705220210LD01	1	217404493	-	3	158848652	+	59	somatic	ASSMB	0.0
C1k_FP1705220210LD01_1:218053493:-_1:218054272:-	FP1705220210LD01	1	218053493	-	1	218054272	-	67	somatic	ASDIS	1.0
C5k_FP1705220210LD01_1:218113670:+_1:218115045:-	FP1705220210LD01	1	218113670	+	1	218115045	-	37	somatic	ASSMB	1.0
C5k_FP1705220210LD01_1:218333114:-_1:218336600:-	FP1705220210LD01	1	218333114	-	1	218336600	-	99	somatic	ASDIS	1.0
C5k_FP1705220210LD01_1:218634576:+_1:218636151:+	FP1705220210LD01	1	218634576	+	1	218636151	+	33	somatic	DSCRD	1.0
Ctran_FP1705220210LD01_1:219985949:-_3:47627829:+	FP1705220210LD01	1	219985949	-	3	47627829	+	53	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_1:221656489:+_5:39794455:+	FP1705220210LD01	1	221656489	+	5	39794455	+	32	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_1:221872646:+_18:10207516:+	FP1705220210LD01	1	221872646	+	18	10207516	+	39	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_1:221873077:-_18:10206991:-	FP1705220210LD01	1	221873077	-	18	10206991	-	67	somatic	ASDIS	0.0
C5k_FP1705220210LD01_1:226017769:+_1:226021132:-	FP1705220210LD01	1	226017769	+	1	226021132	-	10	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_1:226152881:+_6:12092810:-	FP1705220210LD01	1	226152881	+	6	12092810	-	31	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_1:226152887:-_6:12092793:+	FP1705220210LD01	1	226152887	-	6	12092793	+	99	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_1:228009365:+_4:126134593:+	FP1705220210LD01	1	228009365	+	4	126134593	+	22	somatic	DSCRD	0.0
C10k_FP1705220210LD01_1:230843437:+_1:230852803:-	FP1705220210LD01	1	230843437	+	1	230852803	-	33	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_1:234050872:-_3:165830095:+	FP1705220210LD01	1	234050872	-	3	165830095	+	86	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_1:234050877:+_3:165830105:-	FP1705220210LD01	1	234050877	+	3	165830105	-	43	somatic	ASSMB	0.0
C5k_FP1705220210LD01_1:239838272:+_1:239842602:-	FP1705220210LD01	1	239838272	+	1	239842602	-	25	somatic	DSCRD	1.0
C100k_FP1705220210LD01_1:243291743:+_1:243312972:-	FP1705220210LD01	1	243291743	+	1	243312972	-	89	somatic	ASSMB	1.0
C5k_FP1705220210LD01_1:244121840:+_1:244126603:-	FP1705220210LD01	1	244121840	+	1	244126603	-	15	somatic	ASSMB	1.0
C10k_FP1705220210LD01_1:245015880:+_1:245022184:-	FP1705220210LD01	1	245015880	+	1	245022184	-	37	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_1:245098548:-_10:133063522:+	FP1705220210LD01	1	245098548	-	10	133063522	+	16	somatic	ASSMB	0.0
C5k_FP1705220210LD01_1:246808866:+_1:246812135:-	FP1705220210LD01	1	246808866	+	1	246812135	-	15	somatic	DSCRD	1.0
C10k_FP1705220210LD01_1:246816049:+_1:246822868:-	FP1705220210LD01	1	246816049	+	1	246822868	-	32	somatic	ASSMB	1.0
C1k_FP1705220210LD01_1:247881245:+_1:247881695:-	FP1705220210LD01	1	247881245	+	1	247881695	-	32	somatic	ASDIS	1.0
C10k_FP1705220210LD01_2:1046844:+_2:1056809:-	FP1705220210LD01	2	1046844	+	2	1056809	-	54	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_2:2225914:-_15:97701406:-	FP1705220210LD01	2	2225914	-	15	97701406	-	48	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_2:2225969:+_15:97696609:+	FP1705220210LD01	2	2225969	+	15	97696609	+	29	somatic	DSCRD	0.0
C100k_FP1705220210LD01_2:3407161:+_2:3419323:-	FP1705220210LD01	2	3407161	+	2	3419323	-	10	somatic	TSI_L	0.0
Ctran_FP1705220210LD01_2:3407161:+_11:66130001:-	FP1705220210LD01	2	3407161	+	11	66130001	-	54	somatic	TSI_G	0.0
C5k_FP1705220210LD01_2:3407208:-_2:3409438:+	FP1705220210LD01	2	3407208	-	2	3409438	+	20	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_2:3407998:-_11:66130387:+	FP1705220210LD01	2	3407998	-	11	66130387	+	16	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_2:3419463:+_11:66130001:-	FP1705220210LD01	2	3419463	+	11	66130001	-	25	somatic	TSI_L	0.0
C5k_FP1705220210LD01_2:5907178:+_2:5908631:-	FP1705220210LD01	2	5907178	+	2	5908631	-	25	somatic	ASDIS	1.0
C1k_FP1705220210LD01_2:6964236:+_2:6964663:-	FP1705220210LD01	2	6964236	+	2	6964663	-	51	somatic	ASDIS	1.0
C100k_FP1705220210LD01_2:7405978:+_2:7489362:-	FP1705220210LD01	2	7405978	+	2	7489362	-	20	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_2:7820174:-_6:20169002:-	FP1705220210LD01	2	7820174	-	6	20169002	-	15	somatic	DSCRD	0.0
C100k_FP1705220210LD01_2:9189274:+_2:9202112:-	FP1705220210LD01	2	9189274	+	2	9202112	-	20	somatic	ASSMB	1.0
C100k_FP1705220210LD01_2:10118543:-_2:10182756:+	FP1705220210LD01	2	10118543	-	2	10182756	+	10	somatic	DSCRD	1.0
C1k_FP1705220210LD01_2:10366817:+_2:10367357:-	FP1705220210LD01	2	10366817	+	2	10367357	-	11	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:10766934:+_2:10767482:-	FP1705220210LD01	2	10766934	+	2	10767482	-	22	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_2:12293407:+_3:190725700:+	FP1705220210LD01	2	12293407	+	3	190725700	+	14	somatic	DSCRD	0.0
C1k_FP1705220210LD01_2:13861058:+_2:13861780:-	FP1705220210LD01	2	13861058	+	2	13861780	-	16	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_2:14090132:-_22:29066182:+	FP1705220210LD01	2	14090132	-	22	29066182	+	30	somatic	DSCRD	0.0
C100k_FP1705220210LD01_2:20521572:+_2:20539391:-	FP1705220210LD01	2	20521572	+	2	20539391	-	62	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_2:22246330:-_11:71372814:-	FP1705220210LD01	2	22246330	-	11	71372814	-	99	somatic	ASDIS	0.0
C1k_FP1705220210LD01_2:25108116:+_2:25108923:-	FP1705220210LD01	2	25108116	+	2	25108923	-	28	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:26629018:+_2:26629507:-	FP1705220210LD01	2	26629018	+	2	26629507	-	21	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:27443549:+_2:27443904:-	FP1705220210LD01	2	27443549	+	2	27443904	-	40	somatic	ASSMB	1.0
C1M_FP1705220210LD01_2:28624426:-_2:28886632:+	FP1705220210LD01	2	28624426	-	2	28886632	+	26	somatic	ASSMB	1.0
C5k_FP1705220210LD01_2:35488994:+_2:35490586:-	FP1705220210LD01	2	35488994	+	2	35490586	-	66	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:37896173:+_2:37896408:-	FP1705220210LD01	2	37896173	+	2	37896408	-	21	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_2:38709096:-_2:234588695:-	FP1705220210LD01	2	38709096	-	2	234588695	-	82	somatic	ASDIS	0.0
C1k_FP1705220210LD01_2:40882288:+_2:40882575:-	FP1705220210LD01	2	40882288	+	2	40882575	-	32	somatic	ASSMB	1.0
C100k_FP1705220210LD01_2:41655941:+_2:41682912:-	FP1705220210LD01	2	41655941	+	2	41682912	-	55	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_2:48462250:-_8:87715766:-	FP1705220210LD01	2	48462250	-	8	87715766	-	39	somatic	ASDIS	0.0
C1k_FP1705220210LD01_2:51722299:+_2:51722309:-	FP1705220210LD01	2	51722299	+	2	51722309	-	83	somatic	TSI_G	1.0
CBeyond1M_FP1705220210LD01_2:51722299:+_2:54886938:-	FP1705220210LD01	2	51722299	+	2	54886938	-	15	somatic	TSI_L	0.0
CBeyond1M_FP1705220210LD01_2:51722309:-_2:54887412:+	FP1705220210LD01	2	51722309	-	2	54887412	+	47	somatic	TSI_L	0.0
C1k_FP1705220210LD01_2:52005308:+_2:52006168:-	FP1705220210LD01	2	52005308	+	2	52006168	-	26	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_2:55462726:+_12:81532384:-	FP1705220210LD01	2	55462726	+	12	81532384	-	71	somatic	TSI_L	0.0
Ctran_FP1705220210LD01_2:59122813:-_14:59221133:+	FP1705220210LD01	2	59122813	-	14	59221133	+	35	somatic	DSCRD	0.0
C1k_FP1705220210LD01_2:59503535:+_2:59504039:-	FP1705220210LD01	2	59503535	+	2	59504039	-	26	somatic	ASSMB	1.0
C5k_FP1705220210LD01_2:59800506:+_2:59804152:-	FP1705220210LD01	2	59800506	+	2	59804152	-	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:61302667:+_2:61303381:-	FP1705220210LD01	2	61302667	+	2	61303381	-	52	somatic	ASDIS	1.0
C1k_FP1705220210LD01_2:66047127:+_2:66047870:-	FP1705220210LD01	2	66047127	+	2	66047870	-	24	somatic	ASSMB	1.0
C5k_FP1705220210LD01_2:67218625:+_2:67220012:-	FP1705220210LD01	2	67218625	+	2	67220012	-	48	somatic	DSCRD	1.0
C1M_FP1705220210LD01_2:69878895:-_2:70022143:+	FP1705220210LD01	2	69878895	-	2	70022143	+	17	somatic	ASDIS	1.0
C10k_FP1705220210LD01_2:70432558:+_2:70439348:-	FP1705220210LD01	2	70432558	+	2	70439348	-	99	somatic	ASDIS	1.0
C5k_FP1705220210LD01_2:73503269:+_2:73507828:-	FP1705220210LD01	2	73503269	+	2	73507828	-	25	somatic	ASSMB	1.0
C5k_FP1705220210LD01_2:76175195:+_2:76176849:-	FP1705220210LD01	2	76175195	+	2	76176849	-	87	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_2:77572529:-_8:135082457:-	FP1705220210LD01	2	77572529	-	8	135082457	-	50	somatic	DSCRD	0.0
C1k_FP1705220210LD01_2:78140550:+_2:78141311:-	FP1705220210LD01	2	78140550	+	2	78141311	-	29	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_2:78442141:+_2:209707264:-	FP1705220210LD01	2	78442141	+	2	209707264	-	100	somatic	delly_private	0.0
C5k_FP1705220210LD01_2:80420971:+_2:80422044:-	FP1705220210LD01	2	80420971	+	2	80422044	-	31	somatic	ASSMB	1.0
C5k_FP1705220210LD01_2:82343208:+_2:82344573:-	FP1705220210LD01	2	82343208	+	2	82344573	-	52	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_2:95795150:+_6:2785939:+	FP1705220210LD01	2	95795150	+	6	2785939	+	56	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_2:95795174:-_6:2785350:-	FP1705220210LD01	2	95795174	-	6	2785350	-	34	somatic	ASDIS	0.0
C5k_FP1705220210LD01_2:98284342:+_2:98286473:-	FP1705220210LD01	2	98284342	+	2	98286473	-	19	somatic	ASSMB	1.0
C5k_FP1705220210LD01_2:98387996:+_2:98390305:-	FP1705220210LD01	2	98387996	+	2	98390305	-	99	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_2:98465228:-_2:122348078:+	FP1705220210LD01	2	98465228	-	2	122348078	+	62	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_2:103183721:-_7:135887756:-	FP1705220210LD01	2	103183721	-	7	135887756	-	44	somatic	ASDIS	0.0
C1M_FP1705220210LD01_2:103829434:-_2:104757168:+	FP1705220210LD01	2	103829434	-	2	104757168	+	17	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_2:103965556:+_7:125801896:+	FP1705220210LD01	2	103965556	+	7	125801896	+	37	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_2:105256608:-_2:106292628:+	FP1705220210LD01	2	105256608	-	2	106292628	+	23	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_2:107581045:+_2:155646796:-	FP1705220210LD01	2	107581045	+	2	155646796	-	84	somatic	TSI_G	0.0
CBeyond1M_FP1705220210LD01_2:107581115:+_2:178871204:-	FP1705220210LD01	2	107581115	+	2	178871204	-	14	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_2:107591677:-_2:178870980:+	FP1705220210LD01	2	107591677	-	2	178870980	+	92	somatic	TSI_G	0.0
CBeyond1M_FP1705220210LD01_2:107592002:+_2:178871350:-	FP1705220210LD01	2	107592002	+	2	178871350	-	71	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_2:107592166:+_2:155646796:-	FP1705220210LD01	2	107592166	+	2	155646796	-	48	somatic	TSI_L	0.0
CBeyond1M_FP1705220210LD01_2:107592222:-_2:155647067:+	FP1705220210LD01	2	107592222	-	2	155647067	+	63	somatic	ASSMB	0.0
C5k_FP1705220210LD01_2:108595602:+_2:108596747:-	FP1705220210LD01	2	108595602	+	2	108596747	-	99	somatic	ASSMB	1.0
C10k_FP1705220210LD01_2:110423500:+_2:110429864:-	FP1705220210LD01	2	110423500	+	2	110429864	-	83	somatic	DSCRD	1.0
CBeyond1M_FP1705220210LD01_2:110486824:-_2:143174471:-	FP1705220210LD01	2	110486824	-	2	143174471	-	46	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_2:110486835:+_2:143174454:+	FP1705220210LD01	2	110486835	+	2	143174454	+	60	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_2:110931633:+_23:15008032:+	FP1705220210LD01	2	110931633	+	23	15008032	+	99	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_2:110932954:-_23:15007009:-	FP1705220210LD01	2	110932954	-	23	15007009	-	99	somatic	TSI_G	0.0
Ctran_FP1705220210LD01_2:112880415:-_10:83716912:+	FP1705220210LD01	2	112880415	-	10	83716912	+	52	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_2:113752067:-_8:72535184:+	FP1705220210LD01	2	113752067	-	8	72535184	+	28	somatic	TSI_L	0.0
Ctran_FP1705220210LD01_2:113752509:+_8:72534038:+	FP1705220210LD01	2	113752509	+	8	72534038	+	29	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_2:118077384:+_5:39795962:+	FP1705220210LD01	2	118077384	+	5	39795962	+	31	somatic	DSCRD	0.0
C5k_FP1705220210LD01_2:127882439:+_2:127884541:-	FP1705220210LD01	2	127882439	+	2	127884541	-	14	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:130208844:+_2:130209428:-	FP1705220210LD01	2	130208844	+	2	130209428	-	54	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_2:132890395:-_8:135081854:-	FP1705220210LD01	2	132890395	-	8	135081854	-	99	somatic	TSI_G	0.0
C1k_FP1705220210LD01_2:134178887:+_2:134179123:-	FP1705220210LD01	2	134178887	+	2	134179123	-	24	somatic	ASSMB	1.0
C100k_FP1705220210LD01_2:138379839:+_2:138444211:-	FP1705220210LD01	2	138379839	+	2	138444211	-	38	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_2:138917604:+_2:217194437:-	FP1705220210LD01	2	138917604	+	2	217194437	-	56	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_2:138917617:-_2:217194425:+	FP1705220210LD01	2	138917617	-	2	217194425	+	29	somatic	ASSMB	0.0
C1k_FP1705220210LD01_2:139868708:+_2:139869476:-	FP1705220210LD01	2	139868708	+	2	139869476	-	38	somatic	ASSMB	1.0
C1M_FP1705220210LD01_2:140959921:+_2:141144519:-	FP1705220210LD01	2	140959921	+	2	141144519	-	32	somatic	ASSMB	1.0
C1M_FP1705220210LD01_2:141327845:-_2:141681302:+	FP1705220210LD01	2	141327845	-	2	141681302	+	55	somatic	ASSMB	1.0
C10k_FP1705220210LD01_2:141703334:-_2:141710615:+	FP1705220210LD01	2	141703334	-	2	141710615	+	24	somatic	DSCRD	1.0
C1M_FP1705220210LD01_2:141845168:+_2:142058253:-	FP1705220210LD01	2	141845168	+	2	142058253	-	51	somatic	ASSMB	0.0
C1M_FP1705220210LD01_2:141874261:+_2:142070313:-	FP1705220210LD01	2	141874261	+	2	142070313	-	45	somatic	ASSMB	0.0
C5k_FP1705220210LD01_2:142257683:-_2:142260934:+	FP1705220210LD01	2	142257683	-	2	142260934	+	17	somatic	ASSMB	1.0
C100k_FP1705220210LD01_2:142664669:-_2:142691552:+	FP1705220210LD01	2	142664669	-	2	142691552	+	46	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:143342354:+_2:143342798:-	FP1705220210LD01	2	143342354	+	2	143342798	-	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:150843501:+_2:150843827:-	FP1705220210LD01	2	150843501	+	2	150843827	-	11	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:153611984:+_2:153612260:-	FP1705220210LD01	2	153611984	+	2	153612260	-	26	somatic	ASDIS	1.0
C1k_FP1705220210LD01_2:153894874:+_2:153895261:-	FP1705220210LD01	2	153894874	+	2	153895261	-	99	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_2:154002009:-_12:104811258:-	FP1705220210LD01	2	154002009	-	12	104811258	-	15	somatic	DSCRD	0.0
C1k_FP1705220210LD01_2:155646803:+_2:155647061:-	FP1705220210LD01	2	155646803	+	2	155647061	-	19	somatic	TSI_G	1.0
C1k_FP1705220210LD01_2:155647444:+_2:155647699:-	FP1705220210LD01	2	155647444	+	2	155647699	-	33	somatic	TSI_G	1.0
C100k_FP1705220210LD01_2:156596989:+_2:156626754:-	FP1705220210LD01	2	156596989	+	2	156626754	-	59	somatic	ASSMB	1.0
C100k_FP1705220210LD01_2:157968411:+_2:158001099:-	FP1705220210LD01	2	157968411	+	2	158001099	-	40	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_2:164771826:+_9:98465893:+	FP1705220210LD01	2	164771826	+	9	98465893	+	39	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_2:166071976:+_10:82543277:-	FP1705220210LD01	2	166071976	+	10	82543277	-	64	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_2:166074346:-_5:20897817:-	FP1705220210LD01	2	166074346	-	5	20897817	-	24	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_2:166074519:+_9:30762654:-	FP1705220210LD01	2	166074519	+	9	30762654	-	53	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_2:166074573:+_3:138984007:+	FP1705220210LD01	2	166074573	+	3	138984007	+	56	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_2:166075478:-_5:20897906:+	FP1705220210LD01	2	166075478	-	5	20897906	+	30	somatic	DSCRD	0.0
C1k_FP1705220210LD01_2:166075550:+_2:166075996:+	FP1705220210LD01	2	166075550	+	2	166075996	+	27	somatic	DSCRD	1.0
Ctran_FP1705220210LD01_2:166076553:-_4:160351006:+	FP1705220210LD01	2	166076553	-	4	160351006	+	10	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_2:166220461:+_3:55788976:+	FP1705220210LD01	2	166220461	+	3	55788976	+	43	somatic	DSCRD	0.0
C5k_FP1705220210LD01_2:169412430:+_2:169413816:-	FP1705220210LD01	2	169412430	+	2	169413816	-	53	somatic	ASSMB	1.0
C100k_FP1705220210LD01_2:174231917:-_2:174263982:+	FP1705220210LD01	2	174231917	-	2	174263982	+	67	somatic	ASDIS	1.0
C1k_FP1705220210LD01_2:178098449:+_2:178098937:-	FP1705220210LD01	2	178098449	+	2	178098937	-	35	somatic	ASSMB	1.0
C100k_FP1705220210LD01_2:178107014:+_2:178121728:-	FP1705220210LD01	2	178107014	+	2	178121728	-	64	somatic	ASSMB	1.0
C1M_FP1705220210LD01_2:180663216:-_2:180990431:+	FP1705220210LD01	2	180663216	-	2	180990431	+	26	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:181316221:+_2:181317065:-	FP1705220210LD01	2	181316221	+	2	181317065	-	42	somatic	ASSMB	1.0
C100k_FP1705220210LD01_2:182726534:-_2:182772739:+	FP1705220210LD01	2	182726534	-	2	182772739	+	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:184306281:+_2:184306502:-	FP1705220210LD01	2	184306281	+	2	184306502	-	37	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:185834889:-_2:185835332:-	FP1705220210LD01	2	185834889	-	2	185835332	-	96	somatic	ASDIS	1.0
C100k_FP1705220210LD01_2:187405744:-_2:187422803:+	FP1705220210LD01	2	187405744	-	2	187422803	+	21	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_2:196693572:+_4:54368207:-	FP1705220210LD01	2	196693572	+	4	54368207	-	58	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_2:196693792:-_13:25692990:+	FP1705220210LD01	2	196693792	-	13	25692990	+	72	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_2:198367518:-_9:10758487:-	FP1705220210LD01	2	198367518	-	9	10758487	-	46	somatic	TSI_L	0.0
C10k_FP1705220210LD01_2:201533184:+_2:201542764:-	FP1705220210LD01	2	201533184	+	2	201542764	-	32	somatic	ASDIS	1.0
C5k_FP1705220210LD01_2:203173958:+_2:203176569:-	FP1705220210LD01	2	203173958	+	2	203176569	-	24	somatic	DSCRD	1.0
C1k_FP1705220210LD01_2:205007460:+_2:205008180:-	FP1705220210LD01	2	205007460	+	2	205008180	-	19	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_2:207077618:-_11:9771784:-	FP1705220210LD01	2	207077618	-	11	9771784	-	74	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_2:207077703:+_11:9773438:+	FP1705220210LD01	2	207077703	+	11	9773438	+	50	somatic	DSCRD	0.0
C5k_FP1705220210LD01_2:207137379:-_2:207140097:+	FP1705220210LD01	2	207137379	-	2	207140097	+	13	somatic	ASSMB	1.0
C1k_FP1705220210LD01_2:209517994:+_2:209518427:-	FP1705220210LD01	2	209517994	+	2	209518427	-	44	somatic	ASSMB	1.0
C1M_FP1705220210LD01_2:217117023:-_2:217362243:-	FP1705220210LD01	2	217117023	-	2	217362243	-	29	somatic	ASDIS	0.0
C1k_FP1705220210LD01_2:218048681:+_2:218049113:-	FP1705220210LD01	2	218048681	+	2	218049113	-	95	somatic	TSI_G	1.0
Ctran_FP1705220210LD01_2:218048681:+_17:40589618:-	FP1705220210LD01	2	218048681	+	17	40589618	-	65	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_2:218049113:-_17:40589840:+	FP1705220210LD01	2	218049113	-	17	40589840	+	62	somatic	ASSMB	0.0
C5k_FP1705220210LD01_2:232299890:+_2:232301457:-	FP1705220210LD01	2	232299890	+	2	232301457	-	41	somatic	ASDIS	1.0
C1k_FP1705220210LD01_2:234545566:+_2:234546204:-	FP1705220210LD01	2	234545566	+	2	234546204	-	23	somatic	ASSMB	1.0
C100k_FP1705220210LD01_3:215182:-_3:247278:+	FP1705220210LD01	3	215182	-	3	247278	+	99	somatic	DSCRD	1.0
Ctran_FP1705220210LD01_3:1493133:-_13:48244406:-	FP1705220210LD01	3	1493133	-	13	48244406	-	99	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_3:2281324:+_19:48684495:+	FP1705220210LD01	3	2281324	+	19	48684495	+	32	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_3:6008962:-_11:133638804:+	FP1705220210LD01	3	6008962	-	11	133638804	+	59	somatic	ASDIS	0.0
C100k_FP1705220210LD01_3:9114250:+_3:9128153:-	FP1705220210LD01	3	9114250	+	3	9128153	-	29	somatic	DSCRD	1.0
C10k_FP1705220210LD01_3:10253489:+_3:10259073:-	FP1705220210LD01	3	10253489	+	3	10259073	-	13	somatic	ASSMB	1.0
C5k_FP1705220210LD01_3:11396434:+_3:11400858:-	FP1705220210LD01	3	11396434	+	3	11400858	-	47	somatic	ASSMB	1.0
C100k_FP1705220210LD01_3:15366821:-_3:15384869:+	FP1705220210LD01	3	15366821	-	3	15384869	+	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_3:16916519:+_3:16917066:-	FP1705220210LD01	3	16916519	+	3	16917066	-	95	somatic	ASSMB	1.0
C5k_FP1705220210LD01_3:17596369:-_3:17600652:+	FP1705220210LD01	3	17596369	-	3	17600652	+	99	somatic	ASDIS	0.0
C5k_FP1705220210LD01_3:17596487:+_3:17600726:-	FP1705220210LD01	3	17596487	+	3	17600726	-	99	somatic	ASDIS	0.0
C100k_FP1705220210LD01_3:17700829:-_3:17737556:+	FP1705220210LD01	3	17700829	-	3	17737556	+	99	somatic	ASSMB	1.0
C10k_FP1705220210LD01_3:19150713:+_3:19156774:-	FP1705220210LD01	3	19150713	+	3	19156774	-	95	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_3:20586773:-_8:135082731:+	FP1705220210LD01	3	20586773	-	8	135082731	+	17	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_3:32029009:+_13:107870183:-	FP1705220210LD01	3	32029009	+	13	107870183	-	99	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_3:32029016:-_13:107870166:+	FP1705220210LD01	3	32029016	-	13	107870166	+	25	somatic	ASSMB	0.0
C100k_FP1705220210LD01_3:37209543:-_3:37253640:+	FP1705220210LD01	3	37209543	-	3	37253640	+	41	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_3:46260876:+_3:47936135:-	FP1705220210LD01	3	46260876	+	3	47936135	-	59	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_3:49329832:+_16:28048696:-	FP1705220210LD01	3	49329832	+	16	28048696	-	33	somatic	DSCRD	0.0
C1M_FP1705220210LD01_3:50220626:-_3:50834884:+	FP1705220210LD01	3	50220626	-	3	50834884	+	27	somatic	ASSMB	1.0
C1k_FP1705220210LD01_3:52223224:+_3:52223459:-	FP1705220210LD01	3	52223224	+	3	52223459	-	23	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_3:55788662:-_11:24622237:-	FP1705220210LD01	3	55788662	-	11	24622237	-	83	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_3:56424344:-_3:57726265:+	FP1705220210LD01	3	56424344	-	3	57726265	+	42	somatic	ASSMB	1.0
C1k_FP1705220210LD01_3:63022522:+_3:63022840:-	FP1705220210LD01	3	63022522	+	3	63022840	-	68	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_3:63899560:-_13:81737707:+	FP1705220210LD01	3	63899560	-	13	81737707	+	99	somatic	TSI_G	0.0
Ctran_FP1705220210LD01_3:63899560:-_13:81737772:-	FP1705220210LD01	3	63899560	-	13	81737772	-	97	somatic	TSI_L	0.0
C1M_FP1705220210LD01_3:66007986:-_3:66788790:+	FP1705220210LD01	3	66007986	-	3	66788790	+	99	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_3:69460461:-_23:11732777:+	FP1705220210LD01	3	69460461	-	23	11732777	+	80	somatic	DSCRD	0.0
C1M_FP1705220210LD01_3:69481914:+_3:69590305:-	FP1705220210LD01	3	69481914	+	3	69590305	-	99	somatic	ASDIS	1.0
CBeyond1M_FP1705220210LD01_3:69590428:+_3:119927107:-	FP1705220210LD01	3	69590428	+	3	119927107	-	60	somatic	ASSMB	0.0
C1k_FP1705220210LD01_3:74759161:+_3:74759460:-	FP1705220210LD01	3	74759161	+	3	74759460	-	70	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_3:83534197:-_11:7709492:+	FP1705220210LD01	3	83534197	-	11	7709492	+	38	somatic	ASDIS	0.0
C100k_FP1705220210LD01_3:86792293:+_3:86860390:-	FP1705220210LD01	3	86792293	+	3	86860390	-	59	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_3:96519379:+_4:126134740:+	FP1705220210LD01	3	96519379	+	4	126134740	+	25	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_3:96926337:+_3:116940478:-	FP1705220210LD01	3	96926337	+	3	116940478	-	51	somatic	ASSMB	0.0
C1k_FP1705220210LD01_3:104012386:+_3:104012966:-	FP1705220210LD01	3	104012386	+	3	104012966	-	20	somatic	ASSMB	1.0
C5k_FP1705220210LD01_3:104193651:-_3:104195115:+	FP1705220210LD01	3	104193651	-	3	104195115	+	29	somatic	TSI_L	1.0
C1k_FP1705220210LD01_3:104195115:+_3:104195300:-	FP1705220210LD01	3	104195115	+	3	104195300	-	35	somatic	TSI_G	1.0
C1k_FP1705220210LD01_3:104635255:+_3:104635820:-	FP1705220210LD01	3	104635255	+	3	104635820	-	99	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_3:110853111:-_5:71349058:+	FP1705220210LD01	3	110853111	-	5	71349058	+	55	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_3:110853113:+_5:71349064:-	FP1705220210LD01	3	110853113	+	5	71349064	-	55	somatic	ASDIS	0.0
C1M_FP1705220210LD01_3:111287162:-_3:111654716:+	FP1705220210LD01	3	111287162	-	3	111654716	+	55	somatic	ASDIS	0.0
C100k_FP1705220210LD01_3:111573516:+_3:111605223:-	FP1705220210LD01	3	111573516	+	3	111605223	-	49	somatic	DSCRD	1.0
Ctran_FP1705220210LD01_3:122387171:-_10:5399467:+	FP1705220210LD01	3	122387171	-	10	5399467	+	63	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_3:122387574:-_10:5303294:-	FP1705220210LD01	3	122387574	-	10	5303294	-	54	somatic	ASDIS	0.0
C100k_FP1705220210LD01_3:127032566:+_3:127123945:-	FP1705220210LD01	3	127032566	+	3	127123945	-	38	somatic	ASSMB	1.0
C1M_FP1705220210LD01_3:128920977:-_3:129166895:+	FP1705220210LD01	3	128920977	-	3	129166895	+	27	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_3:132721082:-_3:135524024:-	FP1705220210LD01	3	132721082	-	3	135524024	-	96	somatic	ASDIS	0.0
C5k_FP1705220210LD01_3:134760793:+_3:134762400:-	FP1705220210LD01	3	134760793	+	3	134762400	-	15	somatic	ASDIS	1.0
C100k_FP1705220210LD01_3:138970821:+_3:139005697:-	FP1705220210LD01	3	138970821	+	3	139005697	-	29	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_3:140535052:+_2:166077125:+	FP1705220210LD01	3	140535052	+	2	166077125	+	100	somatic	delly_private	0.0
C100k_FP1705220210LD01_3:141745668:+_3:141757264:-	FP1705220210LD01	3	141745668	+	3	141757264	-	29	somatic	ASSMB	1.0
C5k_FP1705220210LD01_3:146488063:+_3:146490113:-	FP1705220210LD01	3	146488063	+	3	146490113	-	21	somatic	ASDIS	1.0
C1k_FP1705220210LD01_3:148864671:+_3:148865039:-	FP1705220210LD01	3	148864671	+	3	148865039	-	39	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_3:149438964:+_6:16147324:-	FP1705220210LD01	3	149438964	+	6	16147324	-	73	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_3:149438977:-_6:16148320:+	FP1705220210LD01	3	149438977	-	6	16148320	+	73	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_3:149958124:-_24:24479473:+	FP1705220210LD01	3	149958124	-	24	24479473	+	38	somatic	ASSMB	0.0
C1k_FP1705220210LD01_3:151623405:-_3:151623714:-	FP1705220210LD01	3	151623405	-	3	151623714	-	44	somatic	ASDIS	1.0
C5k_FP1705220210LD01_3:159553652:-_3:159554990:-	FP1705220210LD01	3	159553652	-	3	159554990	-	99	somatic	TSI_G	0.0
Ctran_FP1705220210LD01_3:159554971:+_10:18742047:-	FP1705220210LD01	3	159554971	+	10	18742047	-	86	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_3:159554990:-_10:18741547:-	FP1705220210LD01	3	159554990	-	10	18741547	-	99	somatic	TSI_L	0.0
Ctran_FP1705220210LD01_3:161970983:+_1:199440237:+	FP1705220210LD01	3	161970983	+	1	199440237	+	100	somatic	delly_private	0.0
C5k_FP1705220210LD01_3:164735365:+_3:164736743:-	FP1705220210LD01	3	164735365	+	3	164736743	-	19	somatic	ASSMB	0.0
C10k_FP1705220210LD01_3:164735877:-_3:164743949:+	FP1705220210LD01	3	164735877	-	3	164743949	+	49	somatic	ASDIS	0.0
C1M_FP1705220210LD01_3:165769231:+_3:166188409:-	FP1705220210LD01	3	165769231	+	3	166188409	-	62	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_3:167774379:-_16:81629104:+	FP1705220210LD01	3	167774379	-	16	81629104	+	46	somatic	DSCRD	0.0
C5k_FP1705220210LD01_3:168167592:+_3:168168980:-	FP1705220210LD01	3	168167592	+	3	168168980	-	75	somatic	ASSMB	1.0
C1k_FP1705220210LD01_3:172045954:+_3:172046171:-	FP1705220210LD01	3	172045954	+	3	172046171	-	29	somatic	ASSMB	1.0
C5k_FP1705220210LD01_3:178231635:+_3:178233463:-	FP1705220210LD01	3	178231635	+	3	178233463	-	59	somatic	ASDIS	1.0
C1k_FP1705220210LD01_3:181501045:+_3:181501524:-	FP1705220210LD01	3	181501045	+	3	181501524	-	49	somatic	ASDIS	1.0
C5k_FP1705220210LD01_3:183181402:+_3:183183446:-	FP1705220210LD01	3	183181402	+	3	183183446	-	92	somatic	DSCRD	1.0
C100k_FP1705220210LD01_3:187654736:+_3:187687036:-	FP1705220210LD01	3	187654736	+	3	187687036	-	83	somatic	ASDIS	1.0
C100k_FP1705220210LD01_3:189349083:+_3:189359219:-	FP1705220210LD01	3	189349083	+	3	189359219	-	38	somatic	ASSMB	1.0
C1k_FP1705220210LD01_3:194674177:+_3:194674977:-	FP1705220210LD01	3	194674177	+	3	194674977	-	41	somatic	ASSMB	1.0
C100k_FP1705220210LD01_3:195034449:-_3:195130466:+	FP1705220210LD01	3	195034449	-	3	195130466	+	99	somatic	ASDIS	1.0
C100k_FP1705220210LD01_3:197007757:+_3:197025689:-	FP1705220210LD01	3	197007757	+	3	197025689	-	18	somatic	ASSMB	1.0
C1M_FP1705220210LD01_4:10747540:-_4:11106888:+	FP1705220210LD01	4	10747540	-	4	11106888	+	39	somatic	ASDIS	1.0
CBeyond1M_FP1705220210LD01_4:14922007:+_4:58849157:+	FP1705220210LD01	4	14922007	+	4	58849157	+	31	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_4:18392225:+_4:126134564:+	FP1705220210LD01	4	18392225	+	4	126134564	+	23	somatic	DSCRD	0.0
C100k_FP1705220210LD01_4:19122429:+_4:19146569:-	FP1705220210LD01	4	19122429	+	4	19146569	-	38	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_4:21167598:+_12:100095952:+	FP1705220210LD01	4	21167598	+	12	100095952	+	65	somatic	DSCRD	0.0
C1k_FP1705220210LD01_4:21440587:+_4:21440848:-	FP1705220210LD01	4	21440587	+	4	21440848	-	44	somatic	ASDIS	1.0
C10k_FP1705220210LD01_4:21526276:+_4:21536110:-	FP1705220210LD01	4	21526276	+	4	21536110	-	38	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_4:28383907:-_11:110016421:-	FP1705220210LD01	4	28383907	-	11	110016421	-	51	somatic	TSI_L	0.0
Ctran_FP1705220210LD01_4:28383975:+_23:105719712:+	FP1705220210LD01	4	28383975	+	23	105719712	+	21	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_4:35960300:+_23:103728505:-	FP1705220210LD01	4	35960300	+	23	103728505	-	32	somatic	DSCRD	0.0
C1k_FP1705220210LD01_4:40402729:+_4:40403013:-	FP1705220210LD01	4	40402729	+	4	40403013	-	45	somatic	ASSMB	1.0
C5k_FP1705220210LD01_4:45133617:-_4:45134693:-	FP1705220210LD01	4	45133617	-	4	45134693	-	20	somatic	ASDIS	1.0
C1k_FP1705220210LD01_4:45140611:-_4:45140709:+	FP1705220210LD01	4	45140611	-	4	45140709	+	31	somatic	TSI_L	1.0
Ctran_FP1705220210LD01_4:45140848:+_12:47304663:-	FP1705220210LD01	4	45140848	+	12	47304663	-	44	somatic	DSCRD	0.0
C5k_FP1705220210LD01_4:52899906:+_4:52900908:-	FP1705220210LD01	4	52899906	+	4	52900908	-	40	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_4:56128934:-_4:57619070:+	FP1705220210LD01	4	56128934	-	4	57619070	+	27	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_4:56491352:-_16:63984748:-	FP1705220210LD01	4	56491352	-	16	63984748	-	52	somatic	ASDIS	0.0
C10k_FP1705220210LD01_4:57281729:+_4:57288821:-	FP1705220210LD01	4	57281729	+	4	57288821	-	50	somatic	ASSMB	1.0
C1k_FP1705220210LD01_4:58599000:+_4:58599531:-	FP1705220210LD01	4	58599000	+	4	58599531	-	20	somatic	ASSMB	1.0
C1k_FP1705220210LD01_4:63207386:+_4:63208342:-	FP1705220210LD01	4	63207386	+	4	63208342	-	98	somatic	ASSMB	1.0
C1k_FP1705220210LD01_4:67805059:+_4:67806033:-	FP1705220210LD01	4	67805059	+	4	67806033	-	99	somatic	ASSMB	1.0
C10k_FP1705220210LD01_4:78447194:-_4:78453470:+	FP1705220210LD01	4	78447194	-	4	78453470	+	42	somatic	ASDIS	1.0
C1M_FP1705220210LD01_4:85484285:-_4:85763310:+	FP1705220210LD01	4	85484285	-	4	85763310	+	48	somatic	ASDIS	1.0
CBeyond1M_FP1705220210LD01_4:86335736:-_4:97875117:-	FP1705220210LD01	4	86335736	-	4	97875117	-	79	somatic	ASDIS	0.0
C1k_FP1705220210LD01_4:89697359:+_4:89697752:-	FP1705220210LD01	4	89697359	+	4	89697752	-	34	somatic	ASDIS	1.0
C100k_FP1705220210LD01_4:91916030:+_4:91939439:-	FP1705220210LD01	4	91916030	+	4	91939439	-	62	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_4:93503016:-_8:73784325:+	FP1705220210LD01	4	93503016	-	8	73784325	+	99	somatic	ASSMB	0.0
C1M_FP1705220210LD01_4:96917745:-_4:97829772:+	FP1705220210LD01	4	96917745	-	4	97829772	+	21	somatic	DSCRD	1.0
C10k_FP1705220210LD01_4:98063286:+_4:98072667:-	FP1705220210LD01	4	98063286	+	4	98072667	-	54	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_4:101754811:-_8:73784588:+	FP1705220210LD01	4	101754811	-	8	73784588	+	46	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_4:101754896:+_8:73783527:-	FP1705220210LD01	4	101754896	+	8	73783527	-	31	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_4:104840224:-_22:29065394:-	FP1705220210LD01	4	104840224	-	22	29065394	-	53	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_4:105699341:+_9:89848131:-	FP1705220210LD01	4	105699341	+	9	89848131	-	52	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_4:105699346:-_9:89848124:+	FP1705220210LD01	4	105699346	-	9	89848124	+	94	somatic	ASSMB	0.0
C1k_FP1705220210LD01_4:108641815:+_4:108642043:-	FP1705220210LD01	4	108641815	+	4	108642043	-	17	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_4:112629029:-_17:60061188:-	FP1705220210LD01	4	112629029	-	17	60061188	-	23	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_4:112629500:+_16:17297810:-	FP1705220210LD01	4	112629500	+	16	17297810	-	38	somatic	ASSMB	0.0
C5k_FP1705220210LD01_4:112630151:-_4:112633135:-	FP1705220210LD01	4	112630151	-	4	112633135	-	64	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_4:112630856:-_8:118735626:+	FP1705220210LD01	4	112630856	-	8	118735626	+	99	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_4:112631174:+_16:17297884:+	FP1705220210LD01	4	112631174	+	16	17297884	+	26	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_4:112631586:+_16:71504598:+	FP1705220210LD01	4	112631586	+	16	71504598	+	74	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_4:124306660:+_23:149006465:-	FP1705220210LD01	4	124306660	+	23	149006465	-	26	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_4:126135132:+_10:96508760:+	FP1705220210LD01	4	126135132	+	10	96508760	+	56	somatic	DSCRD	0.0
C1M_FP1705220210LD01_4:127026112:-_4:127522068:+	FP1705220210LD01	4	127026112	-	4	127522068	+	53	somatic	ASSMB	1.0
C1M_FP1705220210LD01_4:134068440:-_4:134416869:+	FP1705220210LD01	4	134068440	-	4	134416869	+	45	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_4:135038047:+_9:88670345:-	FP1705220210LD01	4	135038047	+	9	88670345	-	10	somatic	ASDIS	0.0
C1k_FP1705220210LD01_4:143540113:+_4:143540294:-	FP1705220210LD01	4	143540113	+	4	143540294	-	86	somatic	ASSMB	1.0
C10k_FP1705220210LD01_4:148495008:+_4:148501432:-	FP1705220210LD01	4	148495008	+	4	148501432	-	78	somatic	ASDIS	1.0
C1k_FP1705220210LD01_4:148929626:-_4:148930528:-	FP1705220210LD01	4	148929626	-	4	148930528	-	23	somatic	ASDIS	1.0
C100k_FP1705220210LD01_4:151519966:+_4:151560651:-	FP1705220210LD01	4	151519966	+	4	151560651	-	89	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_4:157355710:-_8:135082456:-	FP1705220210LD01	4	157355710	-	8	135082456	-	32	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_4:162894835:+_12:117814367:-	FP1705220210LD01	4	162894835	+	12	117814367	-	48	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_4:163267429:+_20:23413451:+	FP1705220210LD01	4	163267429	+	20	23413451	+	58	somatic	TSI_L	0.0
Ctran_FP1705220210LD01_4:164440884:-_16:4790132:-	FP1705220210LD01	4	164440884	-	16	4790132	-	86	somatic	ASDIS	0.0
C100k_FP1705220210LD01_4:168262444:+_4:168281286:-	FP1705220210LD01	4	168262444	+	4	168281286	-	89	somatic	DSCRD	1.0
C100k_FP1705220210LD01_4:176768737:+_4:176782740:-	FP1705220210LD01	4	176768737	+	4	176782740	-	38	somatic	ASSMB	1.0
C1M_FP1705220210LD01_4:181605148:-_4:182599996:+	FP1705220210LD01	4	181605148	-	4	182599996	+	22	somatic	ASDIS	1.0
C5k_FP1705220210LD01_4:183252960:+_4:183254360:-	FP1705220210LD01	4	183252960	+	4	183254360	-	29	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_4:188755977:+_5:44303788:+	FP1705220210LD01	4	188755977	+	5	44303788	+	25	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_4:190590814:+_6:19771419:+	FP1705220210LD01	4	190590814	+	6	19771419	+	32	somatic	DSCRD	0.0
C5k_FP1705220210LD01_5:1106344:+_5:1110000:-	FP1705220210LD01	5	1106344	+	5	1110000	-	89	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_5:1787565:-_10:23745924:+	FP1705220210LD01	5	1787565	-	10	23745924	+	24	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_5:2577165:+_23:46143127:-	FP1705220210LD01	5	2577165	+	23	46143127	-	25	somatic	ASSMB	0.0
C100k_FP1705220210LD01_5:4566303:+_5:4588197:+	FP1705220210LD01	5	4566303	+	5	4588197	+	14	somatic	ASDIS	1.0
C1k_FP1705220210LD01_5:11659109:-_5:11659573:-	FP1705220210LD01	5	11659109	-	5	11659573	-	72	somatic	TSI_L	1.0
C10k_FP1705220210LD01_5:13300162:+_5:13305193:-	FP1705220210LD01	5	13300162	+	5	13305193	-	49	somatic	ASDIS	1.0
C1k_FP1705220210LD01_5:14101139:+_5:14102137:-	FP1705220210LD01	5	14101139	+	5	14102137	-	10	somatic	ASDIS	1.0
C1k_FP1705220210LD01_5:14232882:+_5:14233366:-	FP1705220210LD01	5	14232882	+	5	14233366	-	21	somatic	ASDIS	1.0
C100k_FP1705220210LD01_5:17045689:-_5:17059613:-	FP1705220210LD01	5	17045689	-	5	17059613	-	44	somatic	ASDIS	0.0
C100k_FP1705220210LD01_5:17045912:+_5:17059603:+	FP1705220210LD01	5	17045912	+	5	17059603	+	47	somatic	ASDIS	1.0
C1M_FP1705220210LD01_5:17119082:-_5:17483396:+	FP1705220210LD01	5	17119082	-	5	17483396	+	54	somatic	ASDIS	1.0
C5k_FP1705220210LD01_5:18747735:+_5:18749683:-	FP1705220210LD01	5	18747735	+	5	18749683	-	21	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_5:20582267:+_5:23207211:-	FP1705220210LD01	5	20582267	+	5	23207211	-	24	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_5:22541338:+_22:29065463:+	FP1705220210LD01	5	22541338	+	22	29065463	+	57	somatic	DSCRD	0.0
C1k_FP1705220210LD01_5:23028263:+_5:23028576:-	FP1705220210LD01	5	23028263	+	5	23028576	-	99	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_5:24534731:+_5:32766165:+	FP1705220210LD01	5	24534731	+	5	32766165	+	29	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_5:24534747:-_5:32766172:-	FP1705220210LD01	5	24534747	-	5	32766172	-	54	somatic	ASDIS	0.0
C1k_FP1705220210LD01_5:25554400:+_5:25555286:-	FP1705220210LD01	5	25554400	+	5	25555286	-	20	somatic	ASSMB	1.0
C5k_FP1705220210LD01_5:26144700:+_5:26146269:-	FP1705220210LD01	5	26144700	+	5	26146269	-	12	somatic	ASSMB	1.0
C100k_FP1705220210LD01_5:26273295:-_5:26284139:+	FP1705220210LD01	5	26273295	-	5	26284139	+	19	somatic	ASSMB	1.0
C1k_FP1705220210LD01_5:27405419:+_5:27405703:-	FP1705220210LD01	5	27405419	+	5	27405703	-	99	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_5:28119982:-_23:80876666:-	FP1705220210LD01	5	28119982	-	23	80876666	-	19	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_5:35926299:+_17:21847116:+	FP1705220210LD01	5	35926299	+	17	21847116	+	27	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_5:36318293:-_5:80313467:-	FP1705220210LD01	5	36318293	-	5	80313467	-	35	somatic	TSI_L	0.0
C100k_FP1705220210LD01_5:36854239:+_5:36928256:-	FP1705220210LD01	5	36854239	+	5	36928256	-	35	somatic	ASSMB	1.0
C1M_FP1705220210LD01_5:37090038:+_5:37845173:+	FP1705220210LD01	5	37090038	+	5	37845173	+	58	somatic	ASDIS	0.0
C1M_FP1705220210LD01_5:37090058:-_5:37845178:-	FP1705220210LD01	5	37090058	-	5	37845178	-	49	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_5:39793803:-_23:66518526:-	FP1705220210LD01	5	39793803	-	23	66518526	-	17	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_5:39794680:+_23:66518600:+	FP1705220210LD01	5	39794680	+	23	66518600	+	47	somatic	DSCRD	0.0
C1k_FP1705220210LD01_5:43975853:+_5:43976387:+	FP1705220210LD01	5	43975853	+	5	43976387	+	80	somatic	DSCRD	1.0
Ctran_FP1705220210LD01_5:46105670:+_8:136299029:+	FP1705220210LD01	5	46105670	+	8	136299029	+	26	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_5:50900321:-_22:29066206:+	FP1705220210LD01	5	50900321	-	22	29066206	+	46	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_5:54917717:-_5:130641284:-	FP1705220210LD01	5	54917717	-	5	130641284	-	99	somatic	ASDIS	0.0
C1k_FP1705220210LD01_5:56794208:+_5:56795077:-	FP1705220210LD01	5	56794208	+	5	56795077	-	97	somatic	ASDIS	1.0
C5k_FP1705220210LD01_5:57132759:+_5:57134521:-	FP1705220210LD01	5	57132759	+	5	57134521	-	70	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_5:59409899:-_14:59221135:+	FP1705220210LD01	5	59409899	-	14	59221135	+	61	somatic	DSCRD	0.0
C10k_FP1705220210LD01_5:60701890:+_5:60710090:-	FP1705220210LD01	5	60701890	+	5	60710090	-	29	somatic	ASSMB	1.0
C1k_FP1705220210LD01_5:72598718:+_5:72599472:-	FP1705220210LD01	5	72598718	+	5	72599472	-	46	somatic	ASDIS	1.0
C1M_FP1705220210LD01_5:72634106:-_5:73172915:+	FP1705220210LD01	5	72634106	-	5	73172915	+	60	somatic	ASDIS	0.0
C1k_FP1705220210LD01_5:73124991:+_5:73125510:-	FP1705220210LD01	5	73124991	+	5	73125510	-	26	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_5:74554193:-_17:7816175:+	FP1705220210LD01	5	74554193	-	17	7816175	+	24	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_5:74554202:+_17:7814793:-	FP1705220210LD01	5	74554202	+	17	7814793	-	34	somatic	ASDIS	0.0
C1k_FP1705220210LD01_5:79391953:-_5:79392561:+	FP1705220210LD01	5	79391953	-	5	79392561	+	11	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_5:82059993:+_5:87415450:+	FP1705220210LD01	5	82059993	+	5	87415450	+	38	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_5:84026091:-_16:82113785:-	FP1705220210LD01	5	84026091	-	16	82113785	-	66	somatic	ASDIS	0.0
C1k_FP1705220210LD01_5:84251987:+_5:84252249:-	FP1705220210LD01	5	84251987	+	5	84252249	-	45	somatic	ASSMB	1.0
C1k_FP1705220210LD01_5:84916067:+_5:84917030:-	FP1705220210LD01	5	84916067	+	5	84917030	-	16	somatic	ASSMB	1.0
C1k_FP1705220210LD01_5:100132896:+_5:100133206:-	FP1705220210LD01	5	100132896	+	5	100133206	-	74	somatic	ASDIS	1.0
C100k_FP1705220210LD01_5:100636236:-_5:100646640:+	FP1705220210LD01	5	100636236	-	5	100646640	+	18	somatic	ASDIS	1.0
C1k_FP1705220210LD01_5:106978177:+_5:106978608:-	FP1705220210LD01	5	106978177	+	5	106978608	-	57	somatic	ASDIS	1.0
C10k_FP1705220210LD01_5:120270629:+_5:120279394:-	FP1705220210LD01	5	120270629	+	5	120279394	-	55	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_5:128484926:-_15:52600281:-	FP1705220210LD01	5	128484926	-	15	52600281	-	70	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_5:128485033:+_15:52599479:-	FP1705220210LD01	5	128485033	+	15	52599479	-	32	somatic	DSCRD	0.0
C1M_FP1705220210LD01_5:134067339:-_5:134651887:+	FP1705220210LD01	5	134067339	-	5	134651887	+	53	somatic	ASDIS	1.0
C100k_FP1705220210LD01_5:149403378:-_5:149449506:+	FP1705220210LD01	5	149403378	-	5	149449506	+	14	somatic	DSCRD	1.0
C1k_FP1705220210LD01_5:150158291:+_5:150158768:-	FP1705220210LD01	5	150158291	+	5	150158768	-	18	somatic	ASSMB	1.0
C5k_FP1705220210LD01_5:151527750:+_5:151531523:-	FP1705220210LD01	5	151527750	+	5	151531523	-	61	somatic	ASSMB	1.0
C100k_FP1705220210LD01_5:155106706:-_5:155118639:+	FP1705220210LD01	5	155106706	-	5	155118639	+	40	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_5:163156250:-_9:14152691:-	FP1705220210LD01	5	163156250	-	9	14152691	-	45	somatic	ASDIS	0.0
C1k_FP1705220210LD01_5:173560710:+_5:173561350:-	FP1705220210LD01	5	173560710	+	5	173561350	-	44	somatic	ASSMB	1.0
C5k_FP1705220210LD01_5:176561466:+_5:176566161:-	FP1705220210LD01	5	176561466	+	5	176566161	-	16	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_5:180122155:-_23:65152664:-	FP1705220210LD01	5	180122155	-	23	65152664	-	97	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_5:180122155:-_23:65154756:+	FP1705220210LD01	5	180122155	-	23	65154756	+	99	somatic	TSI_G	0.0
C1M_FP1705220210LD01_6:788191:-_6:1633462:+	FP1705220210LD01	6	788191	-	6	1633462	+	24	somatic	ASSMB	1.0
C1k_FP1705220210LD01_6:13049645:-_6:13050617:-	FP1705220210LD01	6	13049645	-	6	13050617	-	99	somatic	ASDIS	1.0
C1k_FP1705220210LD01_6:13050629:+_6:13051003:-	FP1705220210LD01	6	13050629	+	6	13051003	-	82	somatic	ASSMB	1.0
C100k_FP1705220210LD01_6:13051019:-_6:13062706:-	FP1705220210LD01	6	13051019	-	6	13062706	-	63	somatic	ASDIS	1.0
C100k_FP1705220210LD01_6:15896570:-_6:15978807:-	FP1705220210LD01	6	15896570	-	6	15978807	-	66	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_6:15897427:+_6:123072455:-	FP1705220210LD01	6	15897427	+	6	123072455	-	44	somatic	ASSMB	0.0
C1M_FP1705220210LD01_6:16406932:-_6:16519801:+	FP1705220210LD01	6	16406932	-	6	16519801	+	11	somatic	ASDIS	0.0
C1M_FP1705220210LD01_6:16419788:-_6:16533105:+	FP1705220210LD01	6	16419788	-	6	16533105	+	21	somatic	ASSMB	0.0
C5k_FP1705220210LD01_6:16710981:+_6:16712271:-	FP1705220210LD01	6	16710981	+	6	16712271	-	15	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_6:16821394:+_19:56374264:-	FP1705220210LD01	6	16821394	+	19	56374264	-	51	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_6:18736506:-_8:135082455:-	FP1705220210LD01	6	18736506	-	8	135082455	-	37	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_6:19772250:-_7:53229130:-	FP1705220210LD01	6	19772250	-	7	53229130	-	76	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_6:19835245:-_9:91727631:-	FP1705220210LD01	6	19835245	-	9	91727631	-	82	somatic	ASDIS	0.0
C5k_FP1705220210LD01_6:35359329:+_6:35364261:-	FP1705220210LD01	6	35359329	+	6	35364261	-	10	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_6:38966546:+_11:77320983:-	FP1705220210LD01	6	38966546	+	11	77320983	-	99	somatic	ASSMB	0.0
C1k_FP1705220210LD01_6:38966554:-_6:38967190:-	FP1705220210LD01	6	38966554	-	6	38967190	-	99	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_6:38967475:+_11:77321402:+	FP1705220210LD01	6	38967475	+	11	77321402	+	45	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_6:38968214:+_11:77322086:+	FP1705220210LD01	6	38968214	+	11	77322086	+	35	somatic	DSCRD	0.0
C1k_FP1705220210LD01_6:40765215:+_6:40765476:-	FP1705220210LD01	6	40765215	+	6	40765476	-	15	somatic	ASSMB	1.0
C1k_FP1705220210LD01_6:63074055:+_6:63074655:-	FP1705220210LD01	6	63074055	+	6	63074655	-	30	somatic	ASSMB	1.0
C5k_FP1705220210LD01_6:68011577:+_6:68015275:-	FP1705220210LD01	6	68011577	+	6	68015275	-	78	somatic	ASDIS	1.0
C5k_FP1705220210LD01_6:70349975:+_6:70351107:-	FP1705220210LD01	6	70349975	+	6	70351107	-	29	somatic	ASSMB	1.0
C5k_FP1705220210LD01_6:80498716:+_6:80500124:-	FP1705220210LD01	6	80498716	+	6	80500124	-	47	somatic	ASSMB	1.0
C5k_FP1705220210LD01_6:82256563:+_6:82260747:-	FP1705220210LD01	6	82256563	+	6	82260747	-	90	somatic	ASSMB	1.0
C100k_FP1705220210LD01_6:84754876:-_6:84791436:+	FP1705220210LD01	6	84754876	-	6	84791436	+	17	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_6:92721992:+_6:95994031:+	FP1705220210LD01	6	92721992	+	6	95994031	+	100	somatic	delly_private	0.0
CBeyond1M_FP1705220210LD01_6:92722002:-_6:95994041:-	FP1705220210LD01	6	92722002	-	6	95994041	-	72	somatic	TSI_L	0.0
CBeyond1M_FP1705220210LD01_6:92722166:+_6:95993157:-	FP1705220210LD01	6	92722166	+	6	95993157	-	43	somatic	TSI_L	0.0
CBeyond1M_FP1705220210LD01_6:92722234:-_6:95993289:-	FP1705220210LD01	6	92722234	-	6	95993289	-	99	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_6:95993169:+_15:57215562:-	FP1705220210LD01	6	95993169	+	15	57215562	-	99	somatic	TSI_G	0.0
Ctran_FP1705220210LD01_6:95993294:+_15:57215571:+	FP1705220210LD01	6	95993294	+	15	57215571	+	41	somatic	TSI_L	0.0
Ctran_FP1705220210LD01_6:95994041:-_15:57215571:+	FP1705220210LD01	6	95994041	-	15	57215571	+	99	somatic	TSI_G	0.0
C5k_FP1705220210LD01_6:98358797:+_6:98363337:-	FP1705220210LD01	6	98358797	+	6	98363337	-	52	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_6:101720659:-_12:71020545:+	FP1705220210LD01	6	101720659	-	12	71020545	+	12	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_6:102843553:-_9:105630616:+	FP1705220210LD01	6	102843553	-	9	105630616	+	39	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_6:102844281:+_7:54080823:-	FP1705220210LD01	6	102844281	+	7	54080823	-	15	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_6:102844810:+_9:105630553:-	FP1705220210LD01	6	102844810	+	9	105630553	-	44	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_6:104785582:+_14:59221109:+	FP1705220210LD01	6	104785582	+	14	59221109	+	35	somatic	DSCRD	0.0
C1k_FP1705220210LD01_6:112484074:+_6:112484769:-	FP1705220210LD01	6	112484074	+	6	112484769	-	41	somatic	ASSMB	1.0
C1k_FP1705220210LD01_6:124628476:+_6:124629301:-	FP1705220210LD01	6	124628476	+	6	124629301	-	99	somatic	ASSMB	1.0
C100k_FP1705220210LD01_6:131194869:+_6:131284183:-	FP1705220210LD01	6	131194869	+	6	131284183	-	28	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_6:133136516:-_15:45509356:-	FP1705220210LD01	6	133136516	-	15	45509356	-	53	somatic	ASDIS	0.0
C5k_FP1705220210LD01_6:140861810:+_6:140866640:-	FP1705220210LD01	6	140861810	+	6	140866640	-	99	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_6:161102989:-_8:129406718:+	FP1705220210LD01	6	161102989	-	8	129406718	+	29	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_6:162965819:-_20:57201405:+	FP1705220210LD01	6	162965819	-	20	57201405	+	29	somatic	ASSMB	0.0
C1k_FP1705220210LD01_6:165435830:+_6:165436587:-	FP1705220210LD01	6	165435830	+	6	165436587	-	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_6:169208036:-_6:169208546:-	FP1705220210LD01	6	169208036	-	6	169208546	-	11	somatic	TSI_L	1.0
Ctran_FP1705220210LD01_6:169208553:+_9:119905170:-	FP1705220210LD01	6	169208553	+	9	119905170	-	17	somatic	TSI_L	0.0
C1M_FP1705220210LD01_6:169522672:-_6:170474845:+	FP1705220210LD01	6	169522672	-	6	170474845	+	10	somatic	ASDIS	1.0
C1k_FP1705220210LD01_7:1759925:+_7:1760239:-	FP1705220210LD01	7	1759925	+	7	1760239	-	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_7:9713863:+_7:9714846:-	FP1705220210LD01	7	9713863	+	7	9714846	-	62	somatic	ASSMB	1.0
C1k_FP1705220210LD01_7:10510916:+_7:10511618:-	FP1705220210LD01	7	10510916	+	7	10511618	-	99	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_7:15066518:-_23:11731445:+	FP1705220210LD01	7	15066518	-	23	11731445	+	14	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_7:18453648:+_7:39603039:+	FP1705220210LD01	7	18453648	+	7	39603039	+	47	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_7:18572151:-_9:101544072:+	FP1705220210LD01	7	18572151	-	9	101544072	+	75	somatic	ASDIS	0.0
C5k_FP1705220210LD01_7:18613465:+_7:18616384:-	FP1705220210LD01	7	18613465	+	7	18616384	-	99	somatic	ASDIS	1.0
C5k_FP1705220210LD01_7:21836910:+_7:21838306:-	FP1705220210LD01	7	21836910	+	7	21838306	-	47	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_7:22642533:+_7:102689203:+	FP1705220210LD01	7	22642533	+	7	102689203	+	100	somatic	delly_private	0.0
CBeyond1M_FP1705220210LD01_7:22642567:-_7:102689226:-	FP1705220210LD01	7	22642567	-	7	102689226	-	86	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_7:39603137:-_9:101875285:-	FP1705220210LD01	7	39603137	-	9	101875285	-	94	somatic	ASDIS	0.0
C100k_FP1705220210LD01_7:46693936:+_7:46760733:-	FP1705220210LD01	7	46693936	+	7	46760733	-	21	somatic	ASDIS	1.0
C100k_FP1705220210LD01_7:51027256:+_7:51068295:-	FP1705220210LD01	7	51027256	+	7	51068295	-	73	somatic	ASDIS	1.0
C5k_FP1705220210LD01_7:55492154:+_7:55496139:-	FP1705220210LD01	7	55492154	+	7	55496139	-	33	somatic	ASSMB	1.0
C1k_FP1705220210LD01_7:56072303:+_7:56073066:-	FP1705220210LD01	7	56072303	+	7	56073066	-	16	somatic	ASDIS	1.0
C100k_FP1705220210LD01_7:57396858:+_7:57445024:-	FP1705220210LD01	7	57396858	+	7	57445024	-	16	somatic	ASSMB	1.0
C1k_FP1705220210LD01_7:63894445:+_7:63895008:-	FP1705220210LD01	7	63894445	+	7	63895008	-	50	somatic	ASSMB	1.0
C1M_FP1705220210LD01_7:65348111:-_7:65715456:+	FP1705220210LD01	7	65348111	-	7	65715456	+	21	somatic	DSCRD	0.0
C5k_FP1705220210LD01_7:65542140:+_7:65543344:-	FP1705220210LD01	7	65542140	+	7	65543344	-	27	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_7:66682942:+_13:74831881:-	FP1705220210LD01	7	66682942	+	13	74831881	-	42	somatic	DSCRD	0.0
C100k_FP1705220210LD01_7:69165549:-_7:69228117:+	FP1705220210LD01	7	69165549	-	7	69228117	+	27	somatic	ASSMB	1.0
C5k_FP1705220210LD01_7:71661660:+_7:71663233:-	FP1705220210LD01	7	71661660	+	7	71663233	-	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_7:73807917:+_7:73808363:-	FP1705220210LD01	7	73807917	+	7	73808363	-	56	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_7:77096681:+_8:73785591:+	FP1705220210LD01	7	77096681	+	8	73785591	+	75	somatic	DSCRD	0.0
C1k_FP1705220210LD01_7:83419053:+_7:83419303:-	FP1705220210LD01	7	83419053	+	7	83419303	-	93	somatic	ASSMB	1.0
C5k_FP1705220210LD01_7:88864307:+_7:88866417:-	FP1705220210LD01	7	88864307	+	7	88866417	-	19	somatic	ASDIS	1.0
C5k_FP1705220210LD01_7:90958524:+_7:90961444:-	FP1705220210LD01	7	90958524	+	7	90961444	-	20	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_7:96530433:-_20:26142403:-	FP1705220210LD01	7	96530433	-	20	26142403	-	73	somatic	TSI_L	0.0
C10k_FP1705220210LD01_7:98730017:+_7:98738840:-	FP1705220210LD01	7	98730017	+	7	98738840	-	99	somatic	ASSMB	1.0
C100k_FP1705220210LD01_7:99733235:-_7:99809973:+	FP1705220210LD01	7	99733235	-	7	99809973	+	31	somatic	ASSMB	1.0
C1k_FP1705220210LD01_7:101887306:+_7:101888125:-	FP1705220210LD01	7	101887306	+	7	101888125	-	33	somatic	ASDIS	1.0
C1k_FP1705220210LD01_7:105631215:-_7:105631566:-	FP1705220210LD01	7	105631215	-	7	105631566	-	38	somatic	ASDIS	1.0
C10k_FP1705220210LD01_7:106470218:+_7:106478642:-	FP1705220210LD01	7	106470218	+	7	106478642	-	10	somatic	DSCRD	1.0
C1k_FP1705220210LD01_7:113889054:+_7:113889385:-	FP1705220210LD01	7	113889054	+	7	113889385	-	29	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_7:124453930:+_7:133683624:+	FP1705220210LD01	7	124453930	+	7	133683624	+	72	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_7:124454105:-_7:133683548:-	FP1705220210LD01	7	124454105	-	7	133683548	-	99	somatic	ASDIS	0.0
C5k_FP1705220210LD01_7:125035055:+_7:125036503:-	FP1705220210LD01	7	125035055	+	7	125036503	-	40	somatic	ASSMB	1.0
C5k_FP1705220210LD01_7:135243616:+_7:135245336:-	FP1705220210LD01	7	135243616	+	7	135245336	-	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_7:135481673:+_7:135482386:-	FP1705220210LD01	7	135481673	+	7	135482386	-	29	somatic	ASDIS	1.0
C1k_FP1705220210LD01_7:138007455:+_7:138007895:-	FP1705220210LD01	7	138007455	+	7	138007895	-	99	somatic	ASSMB	1.0
C5k_FP1705220210LD01_7:139647507:+_7:139651769:-	FP1705220210LD01	7	139647507	+	7	139651769	-	26	somatic	ASSMB	1.0
C10k_FP1705220210LD01_7:141659914:-_7:141668454:+	FP1705220210LD01	7	141659914	-	7	141668454	+	77	somatic	ASSMB	1.0
C5k_FP1705220210LD01_7:142136982:+_7:142139788:-	FP1705220210LD01	7	142136982	+	7	142139788	-	36	somatic	ASSMB	1.0
C1k_FP1705220210LD01_7:142513986:-_7:142514592:+	FP1705220210LD01	7	142513986	-	7	142514592	+	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_7:143190432:+_7:143190693:-	FP1705220210LD01	7	143190432	+	7	143190693	-	25	somatic	ASSMB	1.0
C100k_FP1705220210LD01_7:144530909:-_7:144551682:+	FP1705220210LD01	7	144530909	-	7	144551682	+	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_7:145285535:+_7:145285768:-	FP1705220210LD01	7	145285535	+	7	145285768	-	91	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_7:149050287:-_23:150503941:-	FP1705220210LD01	7	149050287	-	23	150503941	-	58	somatic	TSI_G	0.0
Ctran_FP1705220210LD01_7:155819399:-_23:16389104:+	FP1705220210LD01	7	155819399	-	23	16389104	+	91	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_8:5893940:-_15:68045430:-	FP1705220210LD01	8	5893940	-	15	68045430	-	51	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_8:8844814:-_8:17382933:-	FP1705220210LD01	8	8844814	-	8	17382933	-	37	somatic	TSI_L	0.0
CBeyond1M_FP1705220210LD01_8:8845101:+_8:17382631:+	FP1705220210LD01	8	8845101	+	8	17382631	+	66	somatic	TSI_L	1.0
C1k_FP1705220210LD01_8:24367901:+_8:24368449:-	FP1705220210LD01	8	24367901	+	8	24368449	-	35	somatic	ASSMB	1.0
C100k_FP1705220210LD01_8:26959199:+_8:26969291:-	FP1705220210LD01	8	26959199	+	8	26969291	-	32	somatic	ASDIS	1.0
C1M_FP1705220210LD01_8:27463263:-_8:28014576:+	FP1705220210LD01	8	27463263	-	8	28014576	+	30	somatic	ASSMB	0.0
C1k_FP1705220210LD01_8:27892064:-_8:27892722:-	FP1705220210LD01	8	27892064	-	8	27892722	-	34	somatic	ASDIS	1.0
C1k_FP1705220210LD01_8:28884210:+_8:28885070:-	FP1705220210LD01	8	28884210	+	8	28885070	-	15	somatic	ASSMB	1.0
C1k_FP1705220210LD01_8:36370137:+_8:36370459:-	FP1705220210LD01	8	36370137	+	8	36370459	-	44	somatic	ASSMB	1.0
C100k_FP1705220210LD01_8:40255206:-_8:40332986:+	FP1705220210LD01	8	40255206	-	8	40332986	+	23	somatic	ASDIS	1.0
CBeyond1M_FP1705220210LD01_8:41066669:-_8:85415207:+	FP1705220210LD01	8	41066669	-	8	85415207	+	100	somatic	delly_private	0.0
C100k_FP1705220210LD01_8:41770551:+_8:41792745:-	FP1705220210LD01	8	41770551	+	8	41792745	-	30	somatic	ASDIS	1.0
C100k_FP1705220210LD01_8:41967864:+_8:41984236:-	FP1705220210LD01	8	41967864	+	8	41984236	-	60	somatic	ASSMB	1.0
C1k_FP1705220210LD01_8:42500891:+_8:42501528:-	FP1705220210LD01	8	42500891	+	8	42501528	-	29	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_8:51895781:+_14:59221175:+	FP1705220210LD01	8	51895781	+	14	59221175	+	68	somatic	DSCRD	0.0
C1k_FP1705220210LD01_8:52889645:+_8:52890076:-	FP1705220210LD01	8	52889645	+	8	52890076	-	46	somatic	ASDIS	1.0
C1k_FP1705220210LD01_8:53105025:+_8:53105417:-	FP1705220210LD01	8	53105025	+	8	53105417	-	12	somatic	ASSMB	1.0
C1M_FP1705220210LD01_8:53429571:-_8:53610473:+	FP1705220210LD01	8	53429571	-	8	53610473	+	52	somatic	ASSMB	1.0
C10k_FP1705220210LD01_8:54867663:+_8:54873996:-	FP1705220210LD01	8	54867663	+	8	54873996	-	17	somatic	ASSMB	1.0
C1k_FP1705220210LD01_8:55053302:+_8:55053815:-	FP1705220210LD01	8	55053302	+	8	55053815	-	17	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_8:55203197:+_22:29065968:+	FP1705220210LD01	8	55203197	+	22	29065968	+	19	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_8:56908858:+_8:97329042:-	FP1705220210LD01	8	56908858	+	8	97329042	-	49	somatic	ASSMB	0.0
C1k_FP1705220210LD01_8:57539006:-_8:57539727:-	FP1705220210LD01	8	57539006	-	8	57539727	-	99	somatic	ASDIS	1.0
C5k_FP1705220210LD01_8:69124913:+_8:69126170:-	FP1705220210LD01	8	69124913	+	8	69126170	-	42	somatic	ASSMB	1.0
C1M_FP1705220210LD01_8:71104774:+_8:71253698:-	FP1705220210LD01	8	71104774	+	8	71253698	-	32	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_8:73784175:+_9:81554688:-	FP1705220210LD01	8	73784175	+	9	81554688	-	42	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_8:73784191:-_16:51124277:-	FP1705220210LD01	8	73784191	-	16	51124277	-	55	somatic	ASDIS	0.0
C1k_FP1705220210LD01_8:85414874:-_8:85415221:-	FP1705220210LD01	8	85414874	-	8	85415221	-	100	somatic	delly_private	0.0
Ctran_FP1705220210LD01_8:89925188:-_15:86578558:-	FP1705220210LD01	8	89925188	-	15	86578558	-	95	somatic	ASDIS	0.0
C10k_FP1705220210LD01_8:90643909:+_8:90650890:-	FP1705220210LD01	8	90643909	+	8	90650890	-	23	somatic	ASSMB	1.0
C100k_FP1705220210LD01_8:91342261:-_8:91366288:+	FP1705220210LD01	8	91342261	-	8	91366288	+	35	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_8:95340391:+_10:87121581:+	FP1705220210LD01	8	95340391	+	10	87121581	+	36	somatic	DSCRD	0.0
C1M_FP1705220210LD01_8:102264097:-_8:102499582:+	FP1705220210LD01	8	102264097	-	8	102499582	+	58	somatic	ASDIS	1.0
C10k_FP1705220210LD01_8:103233875:+_8:103243844:-	FP1705220210LD01	8	103233875	+	8	103243844	-	39	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_8:104130507:+_19:9042834:-	FP1705220210LD01	8	104130507	+	19	9042834	-	54	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_8:105703911:+_20:62536485:-	FP1705220210LD01	8	105703911	+	20	62536485	-	51	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_8:105703920:-_20:62536459:+	FP1705220210LD01	8	105703920	-	20	62536459	+	60	somatic	ASDIS	0.0
C5k_FP1705220210LD01_8:109070095:+_8:109072953:-	FP1705220210LD01	8	109070095	+	8	109072953	-	31	somatic	ASDIS	1.0
C1M_FP1705220210LD01_8:111314675:-_8:111724847:-	FP1705220210LD01	8	111314675	-	8	111724847	-	58	somatic	TSI_G	0.0
C1k_FP1705220210LD01_8:111351396:+_8:111352332:-	FP1705220210LD01	8	111351396	+	8	111352332	-	20	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_8:112236045:-_11:7710179:-	FP1705220210LD01	8	112236045	-	11	7710179	-	99	somatic	TSI_G	0.0
C1k_FP1705220210LD01_8:112758434:+_8:112759126:-	FP1705220210LD01	8	112758434	+	8	112759126	-	13	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_8:114916146:+_9:98465860:+	FP1705220210LD01	8	114916146	+	9	98465860	+	79	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_8:119429184:+_8:131714791:-	FP1705220210LD01	8	119429184	+	8	131714791	-	25	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_8:119429548:-_8:131715748:+	FP1705220210LD01	8	119429548	-	8	131715748	+	63	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_8:120171994:+_10:123064526:-	FP1705220210LD01	8	120171994	+	10	123064526	-	51	somatic	ASDIS	0.0
C10k_FP1705220210LD01_8:121429126:+_8:121435817:-	FP1705220210LD01	8	121429126	+	8	121435817	-	21	somatic	ASSMB	1.0
C5k_FP1705220210LD01_8:126411089:+_8:126412676:-	FP1705220210LD01	8	126411089	+	8	126412676	-	22	somatic	DSCRD	0.0
C1k_FP1705220210LD01_8:126411999:+_8:126412595:-	FP1705220210LD01	8	126411999	+	8	126412595	-	14	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_8:126514936:-_8:129598218:-	FP1705220210LD01	8	126514936	-	8	129598218	-	99	somatic	ASDIS	0.0
C1M_FP1705220210LD01_8:128166083:-_8:128282097:+	FP1705220210LD01	8	128166083	-	8	128282097	+	61	somatic	ASSMB	0.0
C1M_FP1705220210LD01_8:128212546:-_8:128405543:+	FP1705220210LD01	8	128212546	-	8	128405543	+	99	somatic	ASDIS	0.0
C100k_FP1705220210LD01_8:128775118:-_8:128831717:+	FP1705220210LD01	8	128775118	-	8	128831717	+	39	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_8:129406702:-_14:59221125:+	FP1705220210LD01	8	129406702	-	14	59221125	+	35	somatic	DSCRD	0.0
C5k_FP1705220210LD01_8:129596841:-_8:129599379:+	FP1705220210LD01	8	129596841	-	8	129599379	+	99	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_8:132013503:+_8:145014080:-	FP1705220210LD01	8	132013503	+	8	145014080	-	53	somatic	TSI_L	0.0
CBeyond1M_FP1705220210LD01_8:132013558:+_8:145013210:-	FP1705220210LD01	8	132013558	+	8	145013210	-	19	somatic	DSCRD	0.0
C1k_FP1705220210LD01_8:138697194:+_8:138697545:-	FP1705220210LD01	8	138697194	+	8	138697545	-	38	somatic	ASDIS	1.0
C1k_FP1705220210LD01_8:139497083:+_8:139497741:-	FP1705220210LD01	8	139497083	+	8	139497741	-	13	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_8:139517107:+_8:142289871:+	FP1705220210LD01	8	139517107	+	8	142289871	+	62	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_8:139524629:-_8:142290163:-	FP1705220210LD01	8	139524629	-	8	142290163	-	42	somatic	TSI_G	0.0
C1M_FP1705220210LD01_8:140921330:+_8:141099642:-	FP1705220210LD01	8	140921330	+	8	141099642	-	39	somatic	ASSMB	1.0
C1k_FP1705220210LD01_8:145704612:+_8:145705221:-	FP1705220210LD01	8	145704612	+	8	145705221	-	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_8:146124418:-_8:146124911:+	FP1705220210LD01	8	146124418	-	8	146124911	+	25	somatic	ASDIS	1.0
C5k_FP1705220210LD01_9:1864767:+_9:1867674:-	FP1705220210LD01	9	1864767	+	9	1867674	-	77	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_9:2878293:-_16:26782716:+	FP1705220210LD01	9	2878293	-	16	26782716	+	74	somatic	ASSMB	0.0
C5k_FP1705220210LD01_9:6457822:+_9:6458860:-	FP1705220210LD01	9	6457822	+	9	6458860	-	48	somatic	ASSMB	1.0
C10k_FP1705220210LD01_9:14451686:+_9:14456914:-	FP1705220210LD01	9	14451686	+	9	14456914	-	47	somatic	ASSMB	1.0
C10k_FP1705220210LD01_9:16089462:+_9:16097363:-	FP1705220210LD01	9	16089462	+	9	16097363	-	73	somatic	ASDIS	1.0
C100k_FP1705220210LD01_9:17858733:+_9:17871002:-	FP1705220210LD01	9	17858733	+	9	17871002	-	99	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_9:20055065:+_9:24103665:-	FP1705220210LD01	9	20055065	+	9	24103665	-	99	somatic	ASSMB	1.0
C1M_FP1705220210LD01_9:36100390:-_9:36214459:+	FP1705220210LD01	9	36100390	-	9	36214459	+	44	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_9:76115190:-_18:57070970:-	FP1705220210LD01	9	76115190	-	18	57070970	-	77	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_9:76387905:-_16:83062922:+	FP1705220210LD01	9	76387905	-	16	83062922	+	50	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_9:76387914:+_16:83062934:-	FP1705220210LD01	9	76387914	+	16	83062934	-	36	somatic	ASSMB	0.0
C100k_FP1705220210LD01_9:81355126:-_9:81368695:+	FP1705220210LD01	9	81355126	-	9	81368695	+	57	somatic	ASDIS	1.0
C1k_FP1705220210LD01_9:81661925:+_9:81662912:-	FP1705220210LD01	9	81661925	+	9	81662912	-	22	somatic	ASSMB	1.0
C5k_FP1705220210LD01_9:85399263:+_9:85401689:-	FP1705220210LD01	9	85399263	+	9	85401689	-	99	somatic	ASDIS	1.0
C1k_FP1705220210LD01_9:94994979:+_9:94995924:-	FP1705220210LD01	9	94994979	+	9	94995924	-	99	somatic	ASSMB	1.0
C10k_FP1705220210LD01_9:99915382:+_9:99923806:-	FP1705220210LD01	9	99915382	+	9	99923806	-	54	somatic	ASSMB	1.0
C1k_FP1705220210LD01_9:116946740:+_9:116947046:-	FP1705220210LD01	9	116946740	+	9	116947046	-	14	somatic	ASSMB	1.0
C100k_FP1705220210LD01_9:118793678:+_9:118815941:-	FP1705220210LD01	9	118793678	+	9	118815941	-	55	somatic	ASSMB	1.0
C1k_FP1705220210LD01_9:127948706:+_9:127949245:-	FP1705220210LD01	9	127948706	+	9	127949245	-	27	somatic	ASSMB	1.0
C1k_FP1705220210LD01_9:128048068:+_9:128048674:-	FP1705220210LD01	9	128048068	+	9	128048674	-	80	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_9:129035368:+_9:131598470:+	FP1705220210LD01	9	129035368	+	9	131598470	+	99	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_9:129035374:-_9:130659363:-	FP1705220210LD01	9	129035374	-	9	130659363	-	70	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_9:135627648:-_20:60932731:-	FP1705220210LD01	9	135627648	-	20	60932731	-	56	somatic	ASDIS	0.0
C1k_FP1705220210LD01_10:2440945:+_10:2441889:-	FP1705220210LD01	10	2440945	+	10	2441889	-	46	somatic	ASDIS	1.0
C100k_FP1705220210LD01_10:2730064:-_10:2798130:+	FP1705220210LD01	10	2730064	-	10	2798130	+	18	somatic	ASSMB	1.0
C1k_FP1705220210LD01_10:4095440:+_10:4095692:-	FP1705220210LD01	10	4095440	+	10	4095692	-	17	somatic	ASSMB	1.0
C1k_FP1705220210LD01_10:8062641:+_10:8063540:-	FP1705220210LD01	10	8062641	+	10	8063540	-	44	somatic	ASDIS	1.0
C100k_FP1705220210LD01_10:9148923:+_10:9185137:-	FP1705220210LD01	10	9148923	+	10	9185137	-	58	somatic	ASDIS	1.0
C1k_FP1705220210LD01_10:16163782:+_10:16164232:-	FP1705220210LD01	10	16163782	+	10	16164232	-	32	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_10:18741667:-_3:159554254:-	FP1705220210LD01	10	18741667	-	3	159554254	-	100	somatic	delly_private	0.0
Ctran_FP1705220210LD01_10:18741677:+_3:159553652:-	FP1705220210LD01	10	18741677	+	3	159553652	-	100	somatic	delly_private	0.0
Ctran_FP1705220210LD01_10:18742030:+_3:159554239:+	FP1705220210LD01	10	18742030	+	3	159554239	+	100	somatic	delly_private	0.0
C1k_FP1705220210LD01_10:18774632:+_10:18774978:-	FP1705220210LD01	10	18774632	+	10	18774978	-	48	somatic	ASSMB	1.0
C100k_FP1705220210LD01_10:19593378:+_10:19629296:-	FP1705220210LD01	10	19593378	+	10	19629296	-	71	somatic	ASSMB	1.0
C10k_FP1705220210LD01_10:21369547:-_10:21378011:+	FP1705220210LD01	10	21369547	-	10	21378011	+	39	somatic	ASDIS	1.0
C1M_FP1705220210LD01_10:21407702:-_10:21528034:+	FP1705220210LD01	10	21407702	-	10	21528034	+	32	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_10:27097198:-_10:66522508:+	FP1705220210LD01	10	27097198	-	10	66522508	+	100	somatic	delly_private	0.0
CBeyond1M_FP1705220210LD01_10:27293189:+_10:66522264:+	FP1705220210LD01	10	27293189	+	10	66522264	+	99	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_10:38705327:-_13:96009506:+	FP1705220210LD01	10	38705327	-	13	96009506	+	34	somatic	ASSMB	0.0
C1k_FP1705220210LD01_10:43311726:+_10:43312246:-	FP1705220210LD01	10	43311726	+	10	43312246	-	14	somatic	ASSMB	1.0
C1M_FP1705220210LD01_10:43785237:-_10:44000245:+	FP1705220210LD01	10	43785237	-	10	44000245	+	35	somatic	ASSMB	1.0
C1k_FP1705220210LD01_10:44643173:+_10:44644016:-	FP1705220210LD01	10	44643173	+	10	44644016	-	43	somatic	ASDIS	1.0
C100k_FP1705220210LD01_10:44909921:+_10:44943929:-	FP1705220210LD01	10	44909921	+	10	44943929	-	39	somatic	ASSMB	1.0
C1k_FP1705220210LD01_10:55185394:+_10:55185941:-	FP1705220210LD01	10	55185394	+	10	55185941	-	46	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_10:57920319:+_10:62698690:-	FP1705220210LD01	10	57920319	+	10	62698690	-	72	somatic	ASSMB	1.0
C5k_FP1705220210LD01_10:66222201:+_10:66226794:-	FP1705220210LD01	10	66222201	+	10	66226794	-	89	somatic	ASSMB	1.0
C1k_FP1705220210LD01_10:68539578:+_10:68539877:-	FP1705220210LD01	10	68539578	+	10	68539877	-	24	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_10:71311178:+_10:103927594:+	FP1705220210LD01	10	71311178	+	10	103927594	+	17	somatic	DSCRD	0.0
C1k_FP1705220210LD01_10:74540972:+_10:74541581:-	FP1705220210LD01	10	74540972	+	10	74541581	-	52	somatic	ASSMB	1.0
C100k_FP1705220210LD01_10:79408180:-_10:79418339:+	FP1705220210LD01	10	79408180	-	10	79418339	+	37	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_10:82554195:-_11:7708983:-	FP1705220210LD01	10	82554195	-	11	7708983	-	14	somatic	DSCRD	0.0
C100k_FP1705220210LD01_10:87154527:+_10:87165806:-	FP1705220210LD01	10	87154527	+	10	87165806	-	54	somatic	ASDIS	1.0
C1M_FP1705220210LD01_10:101606033:-_10:102312621:+	FP1705220210LD01	10	101606033	-	10	102312621	+	42	somatic	ASDIS	1.0
C1k_FP1705220210LD01_10:105827062:+_10:105827317:-	FP1705220210LD01	10	105827062	+	10	105827317	-	99	somatic	ASSMB	1.0
C10k_FP1705220210LD01_10:109212939:+_10:109218140:-	FP1705220210LD01	10	109212939	+	10	109218140	-	33	somatic	ASDIS	1.0
C1k_FP1705220210LD01_10:109244736:+_10:109245183:-	FP1705220210LD01	10	109244736	+	10	109245183	-	33	somatic	ASSMB	1.0
C5k_FP1705220210LD01_10:117997672:+_10:117999122:-	FP1705220210LD01	10	117997672	+	10	117999122	-	38	somatic	ASSMB	1.0
C1k_FP1705220210LD01_10:119077254:+_10:119077884:-	FP1705220210LD01	10	119077254	+	10	119077884	-	36	somatic	ASSMB	1.0
C1M_FP1705220210LD01_10:120983245:-_10:121125487:+	FP1705220210LD01	10	120983245	-	10	121125487	+	26	somatic	ASDIS	1.0
C5k_FP1705220210LD01_10:121621523:+_10:121624966:-	FP1705220210LD01	10	121621523	+	10	121624966	-	25	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_10:124073927:-_17:61486494:-	FP1705220210LD01	10	124073927	-	17	61486494	-	52	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_10:124229597:+_17:61676991:+	FP1705220210LD01	10	124229597	+	17	61676991	+	14	somatic	DSCRD	0.0
C5k_FP1705220210LD01_10:125224413:+_10:125226522:-	FP1705220210LD01	10	125224413	+	10	125226522	-	22	somatic	ASSMB	1.0
C10k_FP1705220210LD01_10:129066314:-_10:129073651:+	FP1705220210LD01	10	129066314	-	10	129073651	+	29	somatic	ASDIS	1.0
CBeyond1M_FP1705220210LD01_11:3890694:-_11:88445047:-	FP1705220210LD01	11	3890694	-	11	88445047	-	59	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_11:10164537:+_11:47691845:-	FP1705220210LD01	11	10164537	+	11	47691845	-	48	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_11:11088038:+_11:111642568:-	FP1705220210LD01	11	11088038	+	11	111642568	-	63	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_11:11088048:-_11:111642545:+	FP1705220210LD01	11	11088048	-	11	111642545	+	24	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_11:15668216:-_11:44191865:+	FP1705220210LD01	11	15668216	-	11	44191865	+	51	somatic	ASSMB	0.0
C1k_FP1705220210LD01_11:16722782:+_11:16723051:-	FP1705220210LD01	11	16722782	+	11	16723051	-	64	somatic	ASSMB	1.0
C10k_FP1705220210LD01_11:17123260:+_11:17131935:-	FP1705220210LD01	11	17123260	+	11	17131935	-	39	somatic	ASSMB	1.0
C1k_FP1705220210LD01_11:20084007:+_11:20084439:-	FP1705220210LD01	11	20084007	+	11	20084439	-	44	somatic	ASSMB	1.0
C100k_FP1705220210LD01_11:28032232:-_11:28045222:+	FP1705220210LD01	11	28032232	-	11	28045222	+	55	somatic	ASSMB	1.0
C1M_FP1705220210LD01_11:38385102:-_11:38775629:+	FP1705220210LD01	11	38385102	-	11	38775629	+	53	somatic	ASSMB	0.0
C1k_FP1705220210LD01_11:38629101:+_11:38629716:-	FP1705220210LD01	11	38629101	+	11	38629716	-	14	somatic	ASSMB	1.0
C100k_FP1705220210LD01_11:40002351:-_11:40033491:+	FP1705220210LD01	11	40002351	-	11	40033491	+	14	somatic	ASDIS	1.0
C1k_FP1705220210LD01_11:44999540:+_11:45000238:-	FP1705220210LD01	11	44999540	+	11	45000238	-	23	somatic	ASDIS	1.0
C5k_FP1705220210LD01_11:46537308:+_11:46539285:-	FP1705220210LD01	11	46537308	+	11	46539285	-	45	somatic	DSCRD	1.0
C100k_FP1705220210LD01_11:47707967:-_11:47765130:+	FP1705220210LD01	11	47707967	-	11	47765130	+	17	somatic	DSCRD	1.0
C100k_FP1705220210LD01_11:47975375:-_11:48018713:+	FP1705220210LD01	11	47975375	-	11	48018713	+	39	somatic	ASDIS	1.0
CBeyond1M_FP1705220210LD01_11:55591518:+_11:59266877:-	FP1705220210LD01	11	55591518	+	11	59266877	-	41	somatic	ASSMB	0.0
C1k_FP1705220210LD01_11:58742438:+_11:58742776:-	FP1705220210LD01	11	58742438	+	11	58742776	-	26	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_11:58824710:+_11:74354975:-	FP1705220210LD01	11	58824710	+	11	74354975	-	47	somatic	ASSMB	0.0
C1k_FP1705220210LD01_11:62839653:-_11:62839911:-	FP1705220210LD01	11	62839653	-	11	62839911	-	36	somatic	TSI_L	0.0
CBeyond1M_FP1705220210LD01_11:62839660:+_11:114861877:-	FP1705220210LD01	11	62839660	+	11	114861877	-	57	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_11:62840108:-_11:114862479:-	FP1705220210LD01	11	62840108	-	11	114862479	-	99	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_11:62840118:+_11:114862488:+	FP1705220210LD01	11	62840118	+	11	114862488	+	48	somatic	TSI_L	0.0
C5k_FP1705220210LD01_11:64220209:+_11:64222009:-	FP1705220210LD01	11	64220209	+	11	64222009	-	20	somatic	ASDIS	1.0
C100k_FP1705220210LD01_11:64466571:-_11:64539661:+	FP1705220210LD01	11	64466571	-	11	64539661	+	29	somatic	ASSMB	1.0
C1k_FP1705220210LD01_11:65196000:+_11:65196949:-	FP1705220210LD01	11	65196000	+	11	65196949	-	66	somatic	ASDIS	1.0
C1k_FP1705220210LD01_11:66024393:+_11:66025157:-	FP1705220210LD01	11	66024393	+	11	66025157	-	23	somatic	ASSMB	1.0
C100k_FP1705220210LD01_11:66880789:+_11:66924317:-	FP1705220210LD01	11	66880789	+	11	66924317	-	26	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_11:67996649:+_11:123049813:+	FP1705220210LD01	11	67996649	+	11	123049813	+	30	somatic	ASDIS	0.0
C10k_FP1705220210LD01_11:68253936:+_11:68259912:-	FP1705220210LD01	11	68253936	+	11	68259912	-	66	somatic	ASSMB	1.0
C5k_FP1705220210LD01_11:69995218:-_11:69996290:+	FP1705220210LD01	11	69995218	-	11	69996290	+	11	somatic	ASSMB	1.0
C1M_FP1705220210LD01_11:73616128:-_11:73827819:+	FP1705220210LD01	11	73616128	-	11	73827819	+	22	somatic	ASDIS	1.0
C5k_FP1705220210LD01_11:77127491:+_11:77129245:-	FP1705220210LD01	11	77127491	+	11	77129245	-	30	somatic	ASSMB	1.0
C100k_FP1705220210LD01_11:79136523:-_11:79233682:+	FP1705220210LD01	11	79136523	-	11	79233682	+	66	somatic	ASDIS	1.0
C100k_FP1705220210LD01_11:80248680:-_11:80286931:+	FP1705220210LD01	11	80248680	-	11	80286931	+	66	somatic	TSI_L	1.0
C10k_FP1705220210LD01_11:80286990:+_11:80293781:-	FP1705220210LD01	11	80286990	+	11	80293781	-	25	somatic	DSCRD	1.0
C100k_FP1705220210LD01_11:80418510:-_11:80512952:+	FP1705220210LD01	11	80418510	-	11	80512952	+	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_11:80525765:+_11:80526229:-	FP1705220210LD01	11	80525765	+	11	80526229	-	31	somatic	ASSMB	1.0
C5k_FP1705220210LD01_11:84633534:+_11:84634626:-	FP1705220210LD01	11	84633534	+	11	84634626	-	39	somatic	ASDIS	1.0
C5k_FP1705220210LD01_11:85307818:-_11:85309042:+	FP1705220210LD01	11	85307818	-	11	85309042	+	99	somatic	ASSMB	1.0
C1k_FP1705220210LD01_11:86239284:+_11:86240257:-	FP1705220210LD01	11	86239284	+	11	86240257	-	41	somatic	ASSMB	1.0
C5k_FP1705220210LD01_11:87045136:+_11:87046472:-	FP1705220210LD01	11	87045136	+	11	87046472	-	67	somatic	ASDIS	1.0
C1k_FP1705220210LD01_11:99446635:+_11:99446950:-	FP1705220210LD01	11	99446635	+	11	99446950	-	47	somatic	ASSMB	1.0
C1k_FP1705220210LD01_11:105840944:+_11:105841745:-	FP1705220210LD01	11	105840944	+	11	105841745	-	77	somatic	ASSMB	1.0
C100k_FP1705220210LD01_11:107328742:-_11:107370983:+	FP1705220210LD01	11	107328742	-	11	107370983	+	68	somatic	ASDIS	1.0
C1M_FP1705220210LD01_11:108740468:-_11:109677476:-	FP1705220210LD01	11	108740468	-	11	109677476	-	99	somatic	ASDIS	0.0
C1M_FP1705220210LD01_11:108740579:+_11:109678365:+	FP1705220210LD01	11	108740579	+	11	109678365	+	25	somatic	DSCRD	0.0
C5k_FP1705220210LD01_11:109773156:-_11:109775535:+	FP1705220210LD01	11	109773156	-	11	109775535	+	32	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_11:109773182:+_11:110787275:+	FP1705220210LD01	11	109773182	+	11	110787275	+	32	somatic	DSCRD	0.0
C5k_FP1705220210LD01_11:109774321:+_11:109775528:-	FP1705220210LD01	11	109774321	+	11	109775528	-	57	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_11:109774325:-_11:110787383:+	FP1705220210LD01	11	109774325	-	11	110787383	+	60	somatic	TSI_L	0.0
C10k_FP1705220210LD01_11:118934442:+_11:118940212:-	FP1705220210LD01	11	118934442	+	11	118940212	-	31	somatic	ASSMB	1.0
C10k_FP1705220210LD01_11:126159485:+_11:126165251:-	FP1705220210LD01	11	126159485	+	11	126165251	-	26	somatic	ASSMB	1.0
C1k_FP1705220210LD01_11:126628856:+_11:126629637:-	FP1705220210LD01	11	126628856	+	11	126629637	-	58	somatic	ASDIS	1.0
C1k_FP1705220210LD01_11:127772019:+_11:127772523:-	FP1705220210LD01	11	127772019	+	11	127772523	-	43	somatic	ASSMB	1.0
C1k_FP1705220210LD01_11:131136412:+_11:131136641:-	FP1705220210LD01	11	131136412	+	11	131136641	-	29	somatic	ASSMB	1.0
C1M_FP1705220210LD01_12:470089:-_12:664180:+	FP1705220210LD01	12	470089	-	12	664180	+	44	somatic	DSCRD	1.0
C1k_FP1705220210LD01_12:4495676:+_12:4495981:-	FP1705220210LD01	12	4495676	+	12	4495981	-	99	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_12:6207943:-_12:50156908:+	FP1705220210LD01	12	6207943	-	12	50156908	+	51	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_12:6208029:+_12:50158798:+	FP1705220210LD01	12	6208029	+	12	50158798	+	87	somatic	DSCRD	0.0
C100k_FP1705220210LD01_12:14910731:-_12:14947403:+	FP1705220210LD01	12	14910731	-	12	14947403	+	33	somatic	ASSMB	1.0
C100k_FP1705220210LD01_12:20102747:+_12:20148106:-	FP1705220210LD01	12	20102747	+	12	20148106	-	36	somatic	ASSMB	1.0
C100k_FP1705220210LD01_12:24579448:-_12:24611640:+	FP1705220210LD01	12	24579448	-	12	24611640	+	54	somatic	ASDIS	1.0
C1M_FP1705220210LD01_12:26388908:-_12:27040867:-	FP1705220210LD01	12	26388908	-	12	27040867	-	70	somatic	TSI_L	1.0
C10k_FP1705220210LD01_12:30426451:+_12:30433351:-	FP1705220210LD01	12	30426451	+	12	30433351	-	30	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_12:33323588:-_18:72447119:+	FP1705220210LD01	12	33323588	-	18	72447119	+	39	somatic	DSCRD	0.0
C100k_FP1705220210LD01_12:34147179:+_12:34162028:-	FP1705220210LD01	12	34147179	+	12	34162028	-	69	somatic	ASDIS	1.0
C10k_FP1705220210LD01_12:44651693:-_12:44656839:+	FP1705220210LD01	12	44651693	-	12	44656839	+	31	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_12:46929210:-_12:48025296:+	FP1705220210LD01	12	46929210	-	12	48025296	+	34	somatic	ASSMB	0.0
C1M_FP1705220210LD01_12:50489129:-_12:50598424:+	FP1705220210LD01	12	50489129	-	12	50598424	+	21	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_12:50704908:+_20:53691498:-	FP1705220210LD01	12	50704908	+	20	53691498	-	59	somatic	TSI_G	0.0
C5k_FP1705220210LD01_12:51970010:+_12:51973416:-	FP1705220210LD01	12	51970010	+	12	51973416	-	48	somatic	ASDIS	1.0
C100k_FP1705220210LD01_12:51974226:+_12:51990550:-	FP1705220210LD01	12	51974226	+	12	51990550	-	64	somatic	ASSMB	1.0
C100k_FP1705220210LD01_12:51991846:+_12:52022784:-	FP1705220210LD01	12	51991846	+	12	52022784	-	12	somatic	DSCRD	0.0
C100k_FP1705220210LD01_12:52010952:+_12:52022785:-	FP1705220210LD01	12	52010952	+	12	52022785	-	48	somatic	TSI_L	0.0
CBeyond1M_FP1705220210LD01_12:52939042:-_12:55613646:+	FP1705220210LD01	12	52939042	-	12	55613646	+	55	somatic	ASSMB	1.0
C100k_FP1705220210LD01_12:57755194:-_12:57767413:+	FP1705220210LD01	12	57755194	-	12	57767413	+	38	somatic	ASSMB	1.0
C100k_FP1705220210LD01_12:61715247:+_12:61734052:-	FP1705220210LD01	12	61715247	+	12	61734052	-	51	somatic	ASSMB	1.0
C5k_FP1705220210LD01_12:63315025:+_12:63318661:-	FP1705220210LD01	12	63315025	+	12	63318661	-	38	somatic	ASDIS	1.0
CBeyond1M_FP1705220210LD01_12:71997885:+_12:103855845:-	FP1705220210LD01	12	71997885	+	12	103855845	-	34	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_12:72300468:-_12:122981453:+	FP1705220210LD01	12	72300468	-	12	122981453	+	47	somatic	ASSMB	0.0
C10k_FP1705220210LD01_12:73059960:+_12:73067436:-	FP1705220210LD01	12	73059960	+	12	73067436	-	82	somatic	ASDIS	1.0
C1k_FP1705220210LD01_12:74275222:+_12:74275642:-	FP1705220210LD01	12	74275222	+	12	74275642	-	34	somatic	ASDIS	1.0
C5k_FP1705220210LD01_12:80016886:+_12:80019926:-	FP1705220210LD01	12	80016886	+	12	80019926	-	46	somatic	DSCRD	1.0
C1k_FP1705220210LD01_12:81911175:+_12:81911832:-	FP1705220210LD01	12	81911175	+	12	81911832	-	65	somatic	ASDIS	1.0
C5k_FP1705220210LD01_12:85760640:+_12:85763424:-	FP1705220210LD01	12	85760640	+	12	85763424	-	19	somatic	ASSMB	1.0
C1M_FP1705220210LD01_12:91181209:+_12:91600180:+	FP1705220210LD01	12	91181209	+	12	91600180	+	63	somatic	ASDIS	0.0
C1M_FP1705220210LD01_12:91181227:-_12:91600191:-	FP1705220210LD01	12	91181227	-	12	91600191	-	79	somatic	ASDIS	0.0
C1M_FP1705220210LD01_12:91182023:+_12:91598826:-	FP1705220210LD01	12	91182023	+	12	91598826	-	65	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_12:96960306:+_14:59221162:+	FP1705220210LD01	12	96960306	+	14	59221162	+	21	somatic	DSCRD	0.0
C1k_FP1705220210LD01_12:97658043:+_12:97658847:-	FP1705220210LD01	12	97658043	+	12	97658847	-	41	somatic	ASSMB	1.0
C1M_FP1705220210LD01_12:98497770:-_12:99045158:+	FP1705220210LD01	12	98497770	-	12	99045158	+	42	somatic	DSCRD	0.0
C1M_FP1705220210LD01_12:98784779:-_12:99401682:+	FP1705220210LD01	12	98784779	-	12	99401682	+	25	somatic	ASSMB	0.0
C1M_FP1705220210LD01_12:102733530:-_12:102947637:+	FP1705220210LD01	12	102733530	-	12	102947637	+	31	somatic	ASSMB	1.0
C5k_FP1705220210LD01_12:103565473:+_12:103568447:-	FP1705220210LD01	12	103565473	+	12	103568447	-	74	somatic	ASDIS	1.0
CBeyond1M_FP1705220210LD01_12:103786738:+_12:123623382:-	FP1705220210LD01	12	103786738	+	12	123623382	-	23	somatic	ASSMB	0.0
C1k_FP1705220210LD01_12:119619354:+_12:119619873:-	FP1705220210LD01	12	119619354	+	12	119619873	-	38	somatic	ASDIS	1.0
C1M_FP1705220210LD01_12:122799854:-_12:122969410:+	FP1705220210LD01	12	122799854	-	12	122969410	+	47	somatic	ASSMB	1.0
C10k_FP1705220210LD01_12:123731472:+_12:123737750:+	FP1705220210LD01	12	123731472	+	12	123737750	+	47	somatic	DSCRD	1.0
C5k_FP1705220210LD01_12:125469194:+_12:125474128:-	FP1705220210LD01	12	125469194	+	12	125474128	-	28	somatic	ASSMB	1.0
C100k_FP1705220210LD01_12:127742540:+_12:127780892:-	FP1705220210LD01	12	127742540	+	12	127780892	-	41	somatic	ASSMB	1.0
C1k_FP1705220210LD01_12:130030086:+_12:130030582:-	FP1705220210LD01	12	130030086	+	12	130030582	-	29	somatic	ASDIS	1.0
CBeyond1M_FP1705220210LD01_13:24155672:-_13:31351615:+	FP1705220210LD01	13	24155672	-	13	31351615	+	56	somatic	ASSMB	0.0
Ctran_FP1705220210LD01_13:32550263:+_18:57070978:-	FP1705220210LD01	13	32550263	+	18	57070978	-	50	somatic	DSCRD	0.0
C1k_FP1705220210LD01_13:37446725:+_13:37447165:-	FP1705220210LD01	13	37446725	+	13	37447165	-	40	somatic	ASSMB	1.0
C100k_FP1705220210LD01_13:58327271:+_13:58338782:-	FP1705220210LD01	13	58327271	+	13	58338782	-	63	somatic	ASSMB	1.0
C1k_FP1705220210LD01_13:64248203:+_13:64249011:-	FP1705220210LD01	13	64248203	+	13	64249011	-	39	somatic	ASSMB	1.0
C1k_FP1705220210LD01_13:65108122:+_13:65108569:-	FP1705220210LD01	13	65108122	+	13	65108569	-	99	somatic	ASSMB	1.0
C100k_FP1705220210LD01_13:69215080:+_13:69254460:-	FP1705220210LD01	13	69215080	+	13	69254460	-	68	somatic	ASSMB	1.0
C1M_FP1705220210LD01_13:69445638:-_13:69949904:+	FP1705220210LD01	13	69445638	-	13	69949904	+	35	somatic	ASSMB	1.0
C10k_FP1705220210LD01_13:69965485:-_13:69975148:+	FP1705220210LD01	13	69965485	-	13	69975148	+	99	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_13:71974567:+_13:80856916:-	FP1705220210LD01	13	71974567	+	13	80856916	-	99	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_13:71975087:-_13:80858427:+	FP1705220210LD01	13	71975087	-	13	80858427	+	95	somatic	ASSMB	0.0
CBeyond1M_FP1705220210LD01_13:77495561:+_13:80886200:-	FP1705220210LD01	13	77495561	+	13	80886200	-	99	somatic	ASSMB	0.0
C5k_FP1705220210LD01_13:90673158:+_13:90676301:-	FP1705220210LD01	13	90673158	+	13	90676301	-	99	somatic	ASSMB	1.0
C10k_FP1705220210LD01_13:90724981:-_13:90731157:-	FP1705220210LD01	13	90724981	-	13	90731157	-	13	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_13:91813164:+_14:59220605:-	FP1705220210LD01	13	91813164	+	14	59220605	-	16	somatic	ASSMB	0.0
C5k_FP1705220210LD01_13:99000305:-_13:99002038:-	FP1705220210LD01	13	99000305	-	13	99002038	-	99	somatic	ASDIS	1.0
C1M_FP1705220210LD01_13:104874281:-_13:105472092:+	FP1705220210LD01	13	104874281	-	13	105472092	+	25	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_13:105642336:-_22:36677690:-	FP1705220210LD01	13	105642336	-	22	36677690	-	19	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_13:105642350:+_22:36678624:-	FP1705220210LD01	13	105642350	+	22	36678624	-	46	somatic	TSI_L	0.0
Ctran_FP1705220210LD01_13:105642350:+_22:36680138:-	FP1705220210LD01	13	105642350	+	22	36680138	-	49	somatic	TSI_G	0.0
C10k_FP1705220210LD01_13:107371739:+_13:107379238:-	FP1705220210LD01	13	107371739	+	13	107379238	-	89	somatic	DSCRD	1.0
C100k_FP1705220210LD01_13:109647285:-_13:109682662:+	FP1705220210LD01	13	109647285	-	13	109682662	+	53	somatic	ASDIS	1.0
C100k_FP1705220210LD01_13:110562771:+_13:110574982:-	FP1705220210LD01	13	110562771	+	13	110574982	-	99	somatic	ASSMB	1.0
C5k_FP1705220210LD01_13:113952975:+_13:113954306:-	FP1705220210LD01	13	113952975	+	13	113954306	-	17	somatic	ASSMB	1.0
C5k_FP1705220210LD01_14:23499444:+_14:23500462:-	FP1705220210LD01	14	23499444	+	14	23500462	-	45	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_14:31150680:+_17:49485119:-	FP1705220210LD01	14	31150680	+	17	49485119	-	49	somatic	ASSMB	0.0
C1M_FP1705220210LD01_14:39655959:-_14:39758018:+	FP1705220210LD01	14	39655959	-	14	39758018	+	99	somatic	ASDIS	1.0
C10k_FP1705220210LD01_14:41190379:+_14:41199579:-	FP1705220210LD01	14	41190379	+	14	41199579	-	10	somatic	DSCRD	1.0
C1k_FP1705220210LD01_14:41453811:+_14:41454049:-	FP1705220210LD01	14	41453811	+	14	41454049	-	91	somatic	ASDIS	1.0
C5k_FP1705220210LD01_14:48213542:+_14:48215224:-	FP1705220210LD01	14	48213542	+	14	48215224	-	41	somatic	ASSMB	1.0
C100k_FP1705220210LD01_14:50970570:+_14:50984106:-	FP1705220210LD01	14	50970570	+	14	50984106	-	37	somatic	ASDIS	1.0
C5k_FP1705220210LD01_14:53671385:+_14:53673675:-	FP1705220210LD01	14	53671385	+	14	53673675	-	24	somatic	ASSMB	1.0
C5k_FP1705220210LD01_14:55374607:+_14:55377828:-	FP1705220210LD01	14	55374607	+	14	55377828	-	11	somatic	ASSMB	1.0
C1k_FP1705220210LD01_14:56888625:+_14:56888820:-	FP1705220210LD01	14	56888625	+	14	56888820	-	32	somatic	ASSMB	1.0
C5k_FP1705220210LD01_14:56956904:+_14:56958384:-	FP1705220210LD01	14	56956904	+	14	56958384	-	19	somatic	ASSMB	1.0
C1k_FP1705220210LD01_14:60791378:+_14:60792115:-	FP1705220210LD01	14	60791378	+	14	60792115	-	26	somatic	ASSMB	1.0
C100k_FP1705220210LD01_14:64567322:-_14:64613674:+	FP1705220210LD01	14	64567322	-	14	64613674	+	68	somatic	ASDIS	1.0
C100k_FP1705220210LD01_14:67478120:-_14:67488831:+	FP1705220210LD01	14	67478120	-	14	67488831	+	17	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_14:67605404:-_14:76840672:-	FP1705220210LD01	14	67605404	-	14	76840672	-	23	somatic	ASDIS	0.0
CBeyond1M_FP1705220210LD01_14:68189103:+_14:76828447:+	FP1705220210LD01	14	68189103	+	14	76828447	+	16	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_14:70352364:+_16:24445918:-	FP1705220210LD01	14	70352364	+	16	24445918	-	92	somatic	ASDIS	0.0
C5k_FP1705220210LD01_14:73939020:+_14:73940376:-	FP1705220210LD01	14	73939020	+	14	73940376	-	37	somatic	ASSMB	1.0
C1M_FP1705220210LD01_14:75037699:-_14:75219044:+	FP1705220210LD01	14	75037699	-	14	75219044	+	35	somatic	ASSMB	1.0
C5k_FP1705220210LD01_14:75687867:+_14:75689566:-	FP1705220210LD01	14	75687867	+	14	75689566	-	35	somatic	ASDIS	1.0
C1k_FP1705220210LD01_14:79907527:+_14:79908112:-	FP1705220210LD01	14	79907527	+	14	79908112	-	54	somatic	ASSMB	1.0
C5k_FP1705220210LD01_14:82555638:+_14:82560320:-	FP1705220210LD01	14	82555638	+	14	82560320	-	26	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_14:85651643:+_14:94127300:-	FP1705220210LD01	14	85651643	+	14	94127300	-	35	somatic	ASSMB	0.0
C100k_FP1705220210LD01_14:89044326:-_14:89075610:-	FP1705220210LD01	14	89044326	-	14	89075610	-	22	somatic	DSCRD	0.0
C100k_FP1705220210LD01_14:89044327:-_14:89078086:-	FP1705220210LD01	14	89044327	-	14	89078086	-	99	somatic	TSI_G	0.0
C1k_FP1705220210LD01_14:89077357:+_14:89078093:-	FP1705220210LD01	14	89077357	+	14	89078093	-	13	somatic	DSCRD	0.0
C5k_FP1705220210LD01_14:93135640:+_14:93136831:-	FP1705220210LD01	14	93135640	+	14	93136831	-	44	somatic	ASSMB	1.0
C100k_FP1705220210LD01_14:96755941:-_14:96832451:+	FP1705220210LD01	14	96755941	-	14	96832451	+	48	somatic	ASDIS	1.0
C10k_FP1705220210LD01_14:101279390:+_14:101285822:-	FP1705220210LD01	14	101279390	+	14	101285822	-	52	somatic	ASDIS	1.0
C10k_FP1705220210LD01_14:103020420:+_14:103026720:-	FP1705220210LD01	14	103020420	+	14	103026720	-	29	somatic	ASSMB	1.0
C10k_FP1705220210LD01_14:104386629:+_14:104396258:-	FP1705220210LD01	14	104386629	+	14	104396258	-	40	somatic	ASSMB	1.0
C1M_FP1705220210LD01_14:106092707:+_14:106209402:-	FP1705220210LD01	14	106092707	+	14	106209402	-	26	somatic	DSCRD	1.0
C1M_FP1705220210LD01_15:24496201:+_15:24604746:-	FP1705220210LD01	15	24496201	+	15	24604746	-	17	somatic	DSCRD	1.0
C10k_FP1705220210LD01_15:25176131:-_15:25184263:+	FP1705220210LD01	15	25176131	-	15	25184263	+	62	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_15:25955616:+_15:33197502:-	FP1705220210LD01	15	25955616	+	15	33197502	-	11	somatic	ASSMB	0.0
C5k_FP1705220210LD01_15:31989970:+_15:31991604:-	FP1705220210LD01	15	31989970	+	15	31991604	-	31	somatic	ASDIS	1.0
C5k_FP1705220210LD01_15:33675082:+_15:33676100:-	FP1705220210LD01	15	33675082	+	15	33676100	-	22	somatic	ASSMB	1.0
C1k_FP1705220210LD01_15:40632755:+_15:40633154:-	FP1705220210LD01	15	40632755	+	15	40633154	-	37	somatic	ASDIS	1.0
C1k_FP1705220210LD01_15:52600282:+_15:52601152:+	FP1705220210LD01	15	52600282	+	15	52601152	+	39	somatic	ASDIS	1.0
C1k_FP1705220210LD01_15:53125131:+_15:53125371:-	FP1705220210LD01	15	53125131	+	15	53125371	-	41	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_15:57376654:+_15:80524701:-	FP1705220210LD01	15	57376654	+	15	80524701	-	56	somatic	ASSMB	0.0
C1M_FP1705220210LD01_15:59869406:-_15:59976045:+	FP1705220210LD01	15	59869406	-	15	59976045	+	58	somatic	ASDIS	1.0
C1M_FP1705220210LD01_15:60439552:-_15:60895806:+	FP1705220210LD01	15	60439552	-	15	60895806	+	43	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_15:61102824:-_19:59077272:+	FP1705220210LD01	15	61102824	-	19	59077272	+	22	somatic	DSCRD	0.0
C5k_FP1705220210LD01_15:61493186:+_15:61494446:-	FP1705220210LD01	15	61493186	+	15	61494446	-	32	somatic	ASSMB	1.0
C1k_FP1705220210LD01_15:66537096:+_15:66537553:-	FP1705220210LD01	15	66537096	+	15	66537553	-	35	somatic	ASSMB	1.0
C5k_FP1705220210LD01_15:71816831:+_15:71818442:-	FP1705220210LD01	15	71816831	+	15	71818442	-	51	somatic	ASDIS	1.0
C1k_FP1705220210LD01_15:85567191:+_15:85567634:-	FP1705220210LD01	15	85567191	+	15	85567634	-	86	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_15:90063315:+_22:36677829:+	FP1705220210LD01	15	90063315	+	22	36677829	+	39	somatic	ASDIS	0.0
C5k_FP1705220210LD01_15:94212726:+_15:94214334:-	FP1705220210LD01	15	94212726	+	15	94214334	-	56	somatic	ASDIS	1.0
C5k_FP1705220210LD01_15:94806141:+_15:94808457:-	FP1705220210LD01	15	94806141	+	15	94808457	-	15	somatic	ASSMB	1.0
C5k_FP1705220210LD01_15:98047756:+_15:98049482:-	FP1705220210LD01	15	98047756	+	15	98049482	-	99	somatic	ASSMB	1.0
C100k_FP1705220210LD01_15:98957300:-_15:99019196:+	FP1705220210LD01	15	98957300	-	15	99019196	+	27	somatic	ASSMB	0.0
C5k_FP1705220210LD01_15:98988580:+_15:98989976:-	FP1705220210LD01	15	98988580	+	15	98989976	-	30	somatic	ASSMB	1.0
C100k_FP1705220210LD01_16:338680:-_16:398330:+	FP1705220210LD01	16	338680	-	16	398330	+	57	somatic	ASSMB	1.0
C1k_FP1705220210LD01_16:2740647:+_16:2741170:-	FP1705220210LD01	16	2740647	+	16	2741170	-	19	somatic	ASDIS	1.0
C1M_FP1705220210LD01_16:4978857:-_16:5101012:+	FP1705220210LD01	16	4978857	-	16	5101012	+	36	somatic	DSCRD	1.0
CBeyond1M_FP1705220210LD01_16:11810113:-_16:13813574:-	FP1705220210LD01	16	11810113	-	16	13813574	-	10	somatic	ASDIS	0.0
C10k_FP1705220210LD01_16:13554475:-_16:13559790:+	FP1705220210LD01	16	13554475	-	16	13559790	+	17	somatic	ASSMB	1.0
C1M_FP1705220210LD01_16:14960965:+_16:15876084:+	FP1705220210LD01	16	14960965	+	16	15876084	+	37	somatic	ASDIS	1.0
C100k_FP1705220210LD01_16:17397037:+_16:17426322:-	FP1705220210LD01	16	17397037	+	16	17426322	-	28	somatic	ASSMB	1.0
C1k_FP1705220210LD01_16:25783410:+_16:25783710:-	FP1705220210LD01	16	25783410	+	16	25783710	-	38	somatic	ASSMB	1.0
C5k_FP1705220210LD01_16:29640945:+_16:29641975:-	FP1705220210LD01	16	29640945	+	16	29641975	-	44	somatic	ASDIS	1.0
C5k_FP1705220210LD01_16:33834305:+_16:33836148:-	FP1705220210LD01	16	33834305	+	16	33836148	-	49	somatic	ASSMB	1.0
C100k_FP1705220210LD01_16:34510297:+_16:34535749:-	FP1705220210LD01	16	34510297	+	16	34535749	-	22	somatic	ASDIS	1.0
C100k_FP1705220210LD01_16:47523824:-_16:47535325:+	FP1705220210LD01	16	47523824	-	16	47535325	+	55	somatic	ASDIS	1.0
C5k_FP1705220210LD01_16:52666639:+_16:52667835:-	FP1705220210LD01	16	52666639	+	16	52667835	-	38	somatic	ASDIS	1.0
C5k_FP1705220210LD01_16:57887045:-_16:57888102:-	FP1705220210LD01	16	57887045	-	16	57888102	-	23	somatic	ASDIS	0.0
C100k_FP1705220210LD01_16:57887085:+_16:57897998:+	FP1705220210LD01	16	57887085	+	16	57897998	+	27	somatic	DSCRD	0.0
C1k_FP1705220210LD01_16:60926186:+_16:60926683:-	FP1705220210LD01	16	60926186	+	16	60926683	-	37	somatic	ASSMB	1.0
C1k_FP1705220210LD01_16:61421306:+_16:61421762:-	FP1705220210LD01	16	61421306	+	16	61421762	-	27	somatic	ASSMB	1.0
C1k_FP1705220210LD01_16:70592754:+_16:70593652:-	FP1705220210LD01	16	70592754	+	16	70593652	-	59	somatic	ASDIS	1.0
C5k_FP1705220210LD01_16:72688862:+_16:72690111:-	FP1705220210LD01	16	72688862	+	16	72690111	-	40	somatic	DSCRD	1.0
C10k_FP1705220210LD01_16:74047489:+_16:74054498:-	FP1705220210LD01	16	74047489	+	16	74054498	-	29	somatic	ASSMB	1.0
C1k_FP1705220210LD01_16:78862251:+_16:78862537:-	FP1705220210LD01	16	78862251	+	16	78862537	-	24	somatic	ASSMB	1.0
C1M_FP1705220210LD01_16:81434973:-_16:81549773:+	FP1705220210LD01	16	81434973	-	16	81549773	+	26	somatic	ASDIS	1.0
C1k_FP1705220210LD01_16:81569359:+_16:81569643:-	FP1705220210LD01	16	81569359	+	16	81569643	-	44	somatic	ASSMB	1.0
C100k_FP1705220210LD01_16:87515866:-_16:87542720:+	FP1705220210LD01	16	87515866	-	16	87542720	+	26	somatic	ASSMB	1.0
C5k_FP1705220210LD01_17:4911664:+_17:4914048:-	FP1705220210LD01	17	4911664	+	17	4914048	-	11	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_17:8085801:-_24:15538024:+	FP1705220210LD01	17	8085801	-	24	15538024	+	86	somatic	ASDIS	0.0
C1k_FP1705220210LD01_17:8152598:+_17:8153122:-	FP1705220210LD01	17	8152598	+	17	8153122	-	23	somatic	ASSMB	1.0
C1M_FP1705220210LD01_17:9416656:-_17:9587838:+	FP1705220210LD01	17	9416656	-	17	9587838	+	48	somatic	ASSMB	1.0
C10k_FP1705220210LD01_17:11918588:+_17:11924654:-	FP1705220210LD01	17	11918588	+	17	11924654	-	13	somatic	ASSMB	0.0
C10k_FP1705220210LD01_17:11918602:-_17:11925214:+	FP1705220210LD01	17	11918602	-	17	11925214	+	17	somatic	ASSMB	0.0
C1k_FP1705220210LD01_17:15902858:+_17:15903569:-	FP1705220210LD01	17	15902858	+	17	15903569	-	27	somatic	ASDIS	1.0
C1M_FP1705220210LD01_17:17421457:-_17:18127141:+	FP1705220210LD01	17	17421457	-	17	18127141	+	20	somatic	ASSMB	1.0
C1k_FP1705220210LD01_17:21989610:+_17:21989912:-	FP1705220210LD01	17	21989610	+	17	21989912	-	59	somatic	ASDIS	1.0
C1M_FP1705220210LD01_17:26814714:-_17:27365885:+	FP1705220210LD01	17	26814714	-	17	27365885	+	49	somatic	ASSMB	1.0
C100k_FP1705220210LD01_17:27614673:-_17:27706181:+	FP1705220210LD01	17	27614673	-	17	27706181	+	50	somatic	ASSMB	1.0
C1k_FP1705220210LD01_17:28072635:+_17:28072986:-	FP1705220210LD01	17	28072635	+	17	28072986	-	26	somatic	ASDIS	1.0
C1M_FP1705220210LD01_17:39920306:-_17:40034541:+	FP1705220210LD01	17	39920306	-	17	40034541	+	50	somatic	ASSMB	1.0
C1k_FP1705220210LD01_17:41663741:+_17:41664160:-	FP1705220210LD01	17	41663741	+	17	41664160	-	38	somatic	ASDIS	1.0
C10k_FP1705220210LD01_17:50465118:+_17:50470486:-	FP1705220210LD01	17	50465118	+	17	50470486	-	25	somatic	ASSMB	1.0
C1M_FP1705220210LD01_17:58012046:-_17:58349387:+	FP1705220210LD01	17	58012046	-	17	58349387	+	42	somatic	ASSMB	1.0
C1M_FP1705220210LD01_17:59574729:-_17:59709583:+	FP1705220210LD01	17	59574729	-	17	59709583	+	32	somatic	ASSMB	1.0
C1M_FP1705220210LD01_17:63029936:-_17:63194201:+	FP1705220210LD01	17	63029936	-	17	63194201	+	14	somatic	ASSMB	1.0
C5k_FP1705220210LD01_17:64287936:+_17:64292021:-	FP1705220210LD01	17	64287936	+	17	64292021	-	17	somatic	ASSMB	1.0
C100k_FP1705220210LD01_17:79433578:+_17:79445800:-	FP1705220210LD01	17	79433578	+	17	79445800	-	49	somatic	ASSMB	1.0
C10k_FP1705220210LD01_17:79785252:+_17:79793662:-	FP1705220210LD01	17	79785252	+	17	79793662	-	23	somatic	DSCRD	1.0
C1M_FP1705220210LD01_17:80372792:-_17:80530664:+	FP1705220210LD01	17	80372792	-	17	80530664	+	29	somatic	ASSMB	1.0
C1k_FP1705220210LD01_18:691902:+_18:692267:-	FP1705220210LD01	18	691902	+	18	692267	-	28	somatic	ASDIS	1.0
C5k_FP1705220210LD01_18:1340906:+_18:1343767:-	FP1705220210LD01	18	1340906	+	18	1343767	-	50	somatic	ASDIS	1.0
C100k_FP1705220210LD01_18:3557316:-_18:3600179:+	FP1705220210LD01	18	3557316	-	18	3600179	+	44	somatic	ASDIS	1.0
C1k_FP1705220210LD01_18:3965097:+_18:3965645:-	FP1705220210LD01	18	3965097	+	18	3965645	-	55	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_18:12562167:-_18:19469229:+	FP1705220210LD01	18	12562167	-	18	19469229	+	29	somatic	DSCRD	0.0
C1k_FP1705220210LD01_18:14035109:+_18:14035447:-	FP1705220210LD01	18	14035109	+	18	14035447	-	11	somatic	ASSMB	1.0
C5k_FP1705220210LD01_18:22011464:-_18:22014637:+	FP1705220210LD01	18	22011464	-	18	22014637	+	16	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_18:24194279:+_18:29947069:-	FP1705220210LD01	18	24194279	+	18	29947069	-	68	somatic	TSI_L	1.0
C1M_FP1705220210LD01_18:32616947:+_18:33059711:-	FP1705220210LD01	18	32616947	+	18	33059711	-	38	somatic	ASSMB	1.0
C1k_FP1705220210LD01_18:33121738:+_18:33122378:-	FP1705220210LD01	18	33121738	+	18	33122378	-	88	somatic	ASSMB	1.0
C100k_FP1705220210LD01_18:33697146:-_18:33789019:+	FP1705220210LD01	18	33697146	-	18	33789019	+	86	somatic	ASSMB	1.0
C5k_FP1705220210LD01_18:37164892:-_18:37167796:+	FP1705220210LD01	18	37164892	-	18	37167796	+	71	somatic	ASSMB	1.0
C1k_FP1705220210LD01_18:39395667:+_18:39396149:-	FP1705220210LD01	18	39395667	+	18	39396149	-	29	somatic	ASSMB	1.0
C10k_FP1705220210LD01_18:40122065:+_18:40127620:-	FP1705220210LD01	18	40122065	+	18	40127620	-	22	somatic	DSCRD	1.0
C1k_FP1705220210LD01_18:41785491:+_18:41785988:-	FP1705220210LD01	18	41785491	+	18	41785988	-	33	somatic	ASSMB	1.0
C10k_FP1705220210LD01_18:45512771:+_18:45519009:-	FP1705220210LD01	18	45512771	+	18	45519009	-	30	somatic	ASDIS	1.0
C1k_FP1705220210LD01_18:47065612:+_18:47065927:-	FP1705220210LD01	18	47065612	+	18	47065927	-	31	somatic	ASDIS	1.0
C1k_FP1705220210LD01_18:57659228:+_18:57659465:-	FP1705220210LD01	18	57659228	+	18	57659465	-	99	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_18:58165352:-_22:29065963:+	FP1705220210LD01	18	58165352	-	22	29065963	+	13	somatic	DSCRD	0.0
CBeyond1M_FP1705220210LD01_18:58175706:+_18:68914894:-	FP1705220210LD01	18	58175706	+	18	68914894	-	57	somatic	ASSMB	0.0
C1k_FP1705220210LD01_18:67319720:+_18:67320256:-	FP1705220210LD01	18	67319720	+	18	67320256	-	39	somatic	ASSMB	1.0
C5k_FP1705220210LD01_18:71063356:+_18:71065376:-	FP1705220210LD01	18	71063356	+	18	71065376	-	99	somatic	ASSMB	1.0
C10k_FP1705220210LD01_18:77660959:+_18:77667080:-	FP1705220210LD01	18	77660959	+	18	77667080	-	24	somatic	ASSMB	1.0
C10k_FP1705220210LD01_19:1896183:+_19:1902809:-	FP1705220210LD01	19	1896183	+	19	1902809	-	32	somatic	ASSMB	1.0
C5k_FP1705220210LD01_19:2297426:+_19:2298467:-	FP1705220210LD01	19	2297426	+	19	2298467	-	34	somatic	DSCRD	1.0
C5k_FP1705220210LD01_19:6742222:+_19:6744813:-	FP1705220210LD01	19	6742222	+	19	6744813	-	35	somatic	ASSMB	1.0
C5k_FP1705220210LD01_19:7748361:+_19:7753299:+	FP1705220210LD01	19	7748361	+	19	7753299	+	20	somatic	ASDIS	0.0
C1M_FP1705220210LD01_19:7751364:-_19:8251513:-	FP1705220210LD01	19	7751364	-	19	8251513	-	42	somatic	ASDIS	0.0
C100k_FP1705220210LD01_19:15353625:+_19:15383104:-	FP1705220210LD01	19	15353625	+	19	15383104	-	27	somatic	ASSMB	1.0
C5k_FP1705220210LD01_19:16362727:+_19:16365076:-	FP1705220210LD01	19	16362727	+	19	16365076	-	13	somatic	ASDIS	1.0
C5k_FP1705220210LD01_19:19352646:+_19:19355770:-	FP1705220210LD01	19	19352646	+	19	19355770	-	29	somatic	ASSMB	1.0
C100k_FP1705220210LD01_19:19359796:-_19:19454263:+	FP1705220210LD01	19	19359796	-	19	19454263	+	25	somatic	ASDIS	1.0
C100k_FP1705220210LD01_19:36503154:+_19:36543753:-	FP1705220210LD01	19	36503154	+	19	36543753	-	41	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_19:36711658:-_19:39817670:+	FP1705220210LD01	19	36711658	-	19	39817670	+	55	somatic	ASSMB	1.0
C100k_FP1705220210LD01_19:43701018:+_19:43765018:-	FP1705220210LD01	19	43701018	+	19	43765018	-	15	somatic	DSCRD	1.0
C1M_FP1705220210LD01_19:45036386:-_19:45399968:+	FP1705220210LD01	19	45036386	-	19	45399968	+	66	somatic	ASSMB	0.0
C100k_FP1705220210LD01_19:45350613:+_19:45398203:-	FP1705220210LD01	19	45350613	+	19	45398203	-	27	somatic	ASSMB	1.0
C1k_FP1705220210LD01_19:47445669:+_19:47446601:-	FP1705220210LD01	19	47445669	+	19	47446601	-	25	somatic	ASDIS	1.0
C1M_FP1705220210LD01_19:47506805:-_19:47612138:+	FP1705220210LD01	19	47506805	-	19	47612138	+	28	somatic	ASSMB	1.0
C1k_FP1705220210LD01_19:47809975:+_19:47810246:-	FP1705220210LD01	19	47809975	+	19	47810246	-	17	somatic	ASSMB	1.0
C1k_FP1705220210LD01_19:48948123:+_19:48948531:-	FP1705220210LD01	19	48948123	+	19	48948531	-	42	somatic	TSI_L	1.0
C5k_FP1705220210LD01_19:55395023:+_19:55396766:-	FP1705220210LD01	19	55395023	+	19	55396766	-	27	somatic	DSCRD	1.0
C10k_FP1705220210LD01_19:56735960:+_19:56743141:-	FP1705220210LD01	19	56735960	+	19	56743141	-	38	somatic	ASDIS	1.0
C5k_FP1705220210LD01_20:12112563:+_20:12113734:-	FP1705220210LD01	20	12112563	+	20	12113734	-	14	somatic	ASDIS	1.0
C1M_FP1705220210LD01_20:14504476:+_20:14769832:-	FP1705220210LD01	20	14504476	+	20	14769832	-	41	somatic	ASSMB	1.0
CBeyond1M_FP1705220210LD01_20:17868289:-_20:37795517:+	FP1705220210LD01	20	17868289	-	20	37795517	+	20	somatic	TSI_G	0.0
CBeyond1M_FP1705220210LD01_20:20010920:-_20:29875337:+	FP1705220210LD01	20	20010920	-	20	29875337	+	19	somatic	ASDIS	0.0
C5k_FP1705220210LD01_20:24344625:+_20:24345972:-	FP1705220210LD01	20	24344625	+	20	24345972	-	48	somatic	ASSMB	1.0
C5k_FP1705220210LD01_20:25316545:+_20:25318126:-	FP1705220210LD01	20	25316545	+	20	25318126	-	13	somatic	DSCRD	1.0
C1k_FP1705220210LD01_20:29955414:+_20:29955903:-	FP1705220210LD01	20	29955414	+	20	29955903	-	27	somatic	ASDIS	1.0
C1k_FP1705220210LD01_20:33118586:+_20:33119394:-	FP1705220210LD01	20	33118586	+	20	33119394	-	90	somatic	ASSMB	1.0
C5k_FP1705220210LD01_20:33968141:+_20:33972597:-	FP1705220210LD01	20	33968141	+	20	33972597	-	48	somatic	ASSMB	1.0
C1M_FP1705220210LD01_20:34528764:-_20:34804505:+	FP1705220210LD01	20	34528764	-	20	34804505	+	10	somatic	ASSMB	1.0
C10k_FP1705220210LD01_20:37508891:+_20:37515684:-	FP1705220210LD01	20	37508891	+	20	37515684	-	48	somatic	ASSMB	1.0
C5k_FP1705220210LD01_20:39521120:+_20:39523442:-	FP1705220210LD01	20	39521120	+	20	39523442	-	14	somatic	ASSMB	1.0
C1M_FP1705220210LD01_20:44351228:-_20:44540658:+	FP1705220210LD01	20	44351228	-	20	44540658	+	10	somatic	ASSMB	1.0
C1k_FP1705220210LD01_20:57152470:+_20:57152688:-	FP1705220210LD01	20	57152470	+	20	57152688	-	74	somatic	ASSMB	1.0
C1k_FP1705220210LD01_20:59808468:+_20:59809241:-	FP1705220210LD01	20	59808468	+	20	59809241	-	15	somatic	ASDIS	1.0
C10k_FP1705220210LD01_20:62215839:+_20:62225392:-	FP1705220210LD01	20	62215839	+	20	62225392	-	27	somatic	ASDIS	1.0
C1k_FP1705220210LD01_21:44508268:+_21:44508847:-	FP1705220210LD01	21	44508268	+	21	44508847	-	29	somatic	ASSMB	1.0
C5k_FP1705220210LD01_22:17329316:+_22:17330434:-	FP1705220210LD01	22	17329316	+	22	17330434	-	34	somatic	ASSMB	1.0
C100k_FP1705220210LD01_22:30325562:+_22:30351582:-	FP1705220210LD01	22	30325562	+	22	30351582	-	90	somatic	ASSMB	1.0
C5k_FP1705220210LD01_22:36479701:+_22:36482791:-	FP1705220210LD01	22	36479701	+	22	36482791	-	15	somatic	ASSMB	1.0
C5k_FP1705220210LD01_22:37090392:+_22:37091819:-	FP1705220210LD01	22	37090392	+	22	37091819	-	32	somatic	ASSMB	1.0
C5k_FP1705220210LD01_22:37668840:+_22:37670612:-	FP1705220210LD01	22	37668840	+	22	37670612	-	20	somatic	ASDIS	1.0
C10k_FP1705220210LD01_22:40740365:+_22:40747939:-	FP1705220210LD01	22	40740365	+	22	40747939	-	33	somatic	ASSMB	1.0
C100k_FP1705220210LD01_22:41739186:-_22:41808085:+	FP1705220210LD01	22	41739186	-	22	41808085	+	20	somatic	ASSMB	0.0
C1k_FP1705220210LD01_22:41740005:+_22:41740693:+	FP1705220210LD01	22	41740005	+	22	41740693	+	16	somatic	ASDIS	0.0
C1k_FP1705220210LD01_22:42165890:+_22:42166352:-	FP1705220210LD01	22	42165890	+	22	42166352	-	14	somatic	ASSMB	1.0
C1k_FP1705220210LD01_22:42210113:+_22:42210633:-	FP1705220210LD01	22	42210113	+	22	42210633	-	10	somatic	ASSMB	1.0
C1k_FP1705220210LD01_22:43102130:+_22:43102537:-	FP1705220210LD01	22	43102130	+	22	43102537	-	22	somatic	ASDIS	1.0
C5k_FP1705220210LD01_22:46384768:+_22:46387569:-	FP1705220210LD01	22	46384768	+	22	46387569	-	99	somatic	ASDIS	1.0
C1k_FP1705220210LD01_22:46986162:+_22:46986934:-	FP1705220210LD01	22	46986162	+	22	46986934	-	35	somatic	ASDIS	1.0
C100k_FP1705220210LD01_22:47871739:+_22:47909545:-	FP1705220210LD01	22	47871739	+	22	47909545	-	18	somatic	ASSMB	1.0
C5k_FP1705220210LD01_23:2737752:+_23:2738889:-	FP1705220210LD01	23	2737752	+	23	2738889	-	45	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_23:5657428:+_8:135082456:-	FP1705220210LD01	23	5657428	+	8	135082456	-	12	somatic	DSCRD	0.0
C1M_FP1705220210LD01_23:10403091:+_23:10576066:-	FP1705220210LD01	23	10403091	+	23	10576066	-	66	somatic	ASDIS	1.0
C5k_FP1705220210LD01_23:16387458:+_23:16389095:-	FP1705220210LD01	23	16387458	+	23	16389095	-	99	somatic	TSI_G	1.0
C5k_FP1705220210LD01_23:19738565:+_23:19743290:-	FP1705220210LD01	23	19738565	+	23	19743290	-	14	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_23:23578772:-_8:73783527:-	FP1705220210LD01	23	23578772	-	8	73783527	-	24	somatic	DSCRD	0.0
Ctran_FP1705220210LD01_23:23578784:+_8:73784650:+	FP1705220210LD01	23	23578784	+	8	73784650	+	67	somatic	ASDIS	0.0
C1k_FP1705220210LD01_23:25747238:+_23:25747514:-	FP1705220210LD01	23	25747238	+	23	25747514	-	35	somatic	ASSMB	1.0
C5k_FP1705220210LD01_23:28770571:+_23:28772644:-	FP1705220210LD01	23	28770571	+	23	28772644	-	72	somatic	ASDIS	1.0
C5k_FP1705220210LD01_23:30624720:+_23:30629236:-	FP1705220210LD01	23	30624720	+	23	30629236	-	46	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_23:37532252:-_24:18001188:+	FP1705220210LD01	23	37532252	-	24	18001188	+	93	somatic	ASSMB	0.0
C100k_FP1705220210LD01_23:46762630:-_23:46796604:+	FP1705220210LD01	23	46762630	-	23	46796604	+	65	somatic	ASSMB	1.0
C10k_FP1705220210LD01_23:50441136:+_23:50446637:-	FP1705220210LD01	23	50441136	+	23	50446637	-	25	somatic	ASDIS	1.0
C1k_FP1705220210LD01_23:55919944:+_23:55920317:-	FP1705220210LD01	23	55919944	+	23	55920317	-	66	somatic	ASDIS	1.0
C100k_FP1705220210LD01_23:62754623:-_23:62767803:+	FP1705220210LD01	23	62754623	-	23	62767803	+	50	somatic	ASSMB	1.0
C1k_FP1705220210LD01_23:65104441:+_23:65104687:-	FP1705220210LD01	23	65104441	+	23	65104687	-	34	somatic	ASSMB	1.0
C5k_FP1705220210LD01_23:65151007:+_23:65153417:-	FP1705220210LD01	23	65151007	+	23	65153417	-	44	somatic	ASSMB	0.0
C5k_FP1705220210LD01_23:65153249:+_23:65154803:+	FP1705220210LD01	23	65153249	+	23	65154803	+	42	somatic	DSCRD	0.0
C1M_FP1705220210LD01_23:67505754:-_23:67689736:+	FP1705220210LD01	23	67505754	-	23	67689736	+	10	somatic	ASDIS	1.0
C1M_FP1705220210LD01_23:72908653:-_23:73584471:+	FP1705220210LD01	23	72908653	-	23	73584471	+	27	somatic	ASDIS	1.0
C1M_FP1705220210LD01_23:79059642:-_23:79516635:+	FP1705220210LD01	23	79059642	-	23	79516635	+	22	somatic	ASDIS	1.0
C1k_FP1705220210LD01_23:84600166:+_23:84601065:-	FP1705220210LD01	23	84600166	+	23	84601065	-	60	somatic	ASSMB	1.0
C1M_FP1705220210LD01_23:95347583:-_23:96043612:+	FP1705220210LD01	23	95347583	-	23	96043612	+	23	somatic	ASDIS	1.0
Ctran_FP1705220210LD01_23:103720713:+_4:35959956:-	FP1705220210LD01	23	103720713	+	4	35959956	-	100	somatic	delly_private	0.0
Ctran_FP1705220210LD01_23:110050111:+_6:19771185:+	FP1705220210LD01	23	110050111	+	6	19771185	+	100	somatic	delly_private	0.0
C1k_FP1705220210LD01_23:110198300:+_23:110198630:-	FP1705220210LD01	23	110198300	+	23	110198630	-	51	somatic	ASDIS	1.0
C1k_FP1705220210LD01_23:110509668:+_23:110510308:-	FP1705220210LD01	23	110509668	+	23	110510308	-	58	somatic	ASSMB	1.0
C5k_FP1705220210LD01_23:126000517:+_23:126002534:-	FP1705220210LD01	23	126000517	+	23	126002534	-	56	somatic	ASDIS	1.0
C10k_FP1705220210LD01_23:129403430:+_23:129409166:-	FP1705220210LD01	23	129403430	+	23	129409166	-	49	somatic	DSCRD	1.0
C5k_FP1705220210LD01_23:130284539:+_23:130285787:-	FP1705220210LD01	23	130284539	+	23	130285787	-	48	somatic	DSCRD	1.0
C1k_FP1705220210LD01_23:133650641:+_23:133651515:-	FP1705220210LD01	23	133650641	+	23	133651515	-	41	somatic	DSCRD	1.0
C1k_FP1705220210LD01_23:137353900:+_23:137354131:-	FP1705220210LD01	23	137353900	+	23	137354131	-	24	somatic	ASSMB	1.0
C1k_FP1705220210LD01_23:139947355:+_23:139947596:-	FP1705220210LD01	23	139947355	+	23	139947596	-	24	somatic	ASSMB	1.0
C1M_FP1705220210LD01_23:140974505:-_23:141629717:+	FP1705220210LD01	23	140974505	-	23	141629717	+	23	somatic	ASSMB	1.0
C5k_FP1705220210LD01_23:148154782:+_23:148156148:-	FP1705220210LD01	23	148154782	+	23	148156148	-	36	somatic	ASSMB	1.0
Ctran_FP1705220210LD01_24:4807970:+_22:44316739:+	FP1705220210LD01	24	4807970	+	22	44316739	+	39	somatic	ASDIS	0.0
Ctran_FP1705220210LD01_24:4808015:-_22:44316756:-	FP1705220210LD01	24	4808015	-	22	44316756	-	99	somatic	ASDIS	0.0
C1k_FP1705220210LD01_24:17421916:+_24:17422566:-	FP1705220210LD01	24	17421916	+	24	17422566	-	40	somatic	ASSMB	1.0
C100k_FP1705220210LD01_24:21249766:-_24:21274933:+	FP1705220210LD01	24	21249766	-	24	21274933	+	24	somatic	ASSMB	1.0
